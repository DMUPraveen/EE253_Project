CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 540 30 110 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 D:\Programs\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.209790 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
77
5 4049~
219 892 799 0 2 22
0 4 3
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
5130 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 1903 186 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 1924 233 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.90066e-315 5.26354e-315
0
14 Logic Display~
6 1960 232 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.90066e-315 5.30499e-315
0
14 Logic Display~
6 1942 237 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.90066e-315 5.32571e-315
0
14 Logic Display~
6 2123 452 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44974.7 0
0
14 Logic Display~
6 2122 403 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
44974.7 1
0
14 Logic Display~
6 2121 359 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
44974.7 2
0
14 Logic Display~
6 2109 314 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
44974.7 3
0
7 74LS175
131 2021 353 0 14 29
0 3 5 9 8 7 6 13 61 12
62 11 63 10 64
0
0 0 4832 0
7 74LS175
-24 -51 25 -43
3 U15
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 9 13 12 5 4 15 14 10
11 7 6 2 3 1 9 13 12 5
4 15 14 10 11 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
972 0 0
2
44974.7 4
0
9 Inverter~
13 1759 384 0 2 22
0 15 14
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U14A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3472 0 0
2
44974.7 5
0
7 74LS245
64 1874 420 0 18 37
0 65 66 67 68 16 17 18 19 69
70 71 72 9 8 7 6 14 73
0
0 0 4832 0
7 74LS245
-24 -60 25 -52
3 U13
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
44974.7 6
0
7 74LS245
64 1863 256 0 18 37
0 74 75 76 77 20 21 22 23 78
79 80 81 9 8 7 6 15 82
0
0 0 4832 0
7 74LS245
-24 -60 25 -52
3 U12
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
44974.7 7
0
14 Logic Display~
6 1697 305 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44974.7 8
0
14 Logic Display~
6 1696 265 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
44974.7 9
0
14 Logic Display~
6 1697 189 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
44974.7 10
0
14 Logic Display~
6 1695 146 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
44974.7 11
0
14 NO PushButton~
191 1337 286 0 2 5
0 26 2
0
0 0 4704 0
0
2 S8
-9 -17 5 -9
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9323 0 0
2
44974.7 12
0
14 NO PushButton~
191 1338 322 0 2 5
0 24 2
0
0 0 4704 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
317 0 0
2
44974.7 13
0
14 NO PushButton~
191 1339 203 0 2 5
0 27 2
0
0 0 4704 0
0
2 S6
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3108 0 0
2
44974.7 14
0
14 NO PushButton~
191 1340 167 0 2 5
0 28 2
0
0 0 4704 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4299 0 0
2
44974.7 15
0
7 Ground~
168 1541 27 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
44974.7 16
0
2 +V
167 1457 46 0 1 3
0 25
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
44974.7 17
0
6 74LS73
102 1635 303 0 12 25
0 25 25 26 25 25 25 24 25 22
83 23 84
0
0 0 4832 0
6 74LS73
-21 -51 21 -43
3 U11
-11 -52 10 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
6369 0 0
2
44974.7 18
0
6 74LS73
102 1636 184 0 12 25
0 25 25 28 25 25 25 27 25 20
85 21 86
0
0 0 4832 0
6 74LS73
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
9172 0 0
2
44974.7 19
0
5 4049~
219 272 1033 0 2 22
0 4 29
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
7100 0 0
2
44974.7 20
0
14 NO PushButton~
191 213 1131 0 2 5
0 30 31
0
0 0 4704 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3820 0 0
2
44974.7 21
0
14 Logic Display~
6 813 1277 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
44974.7 22
0
14 Logic Display~
6 812 1190 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
44974.7 23
0
14 Logic Display~
6 815 1093 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
44974.7 24
0
4 4017
219 552 1165 0 14 29
0 29 30 34 32 15 33 34 87 88
89 90 91 92 93
0
0 0 6880 0
4 4017
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
44974.7 25
0
5 4049~
219 278 475 0 2 22
0 5 36
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
3951 0 0
2
44974.7 26
0
14 NO PushButton~
191 229 871 0 2 5
0 38 31
0
0 0 4704 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8885 0 0
2
44974.7 27
0
5 4049~
219 229 527 0 2 22
0 38 39
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
3780 0 0
2
44974.7 28
0
9 2-In AND~
219 240 567 0 3 22
0 39 41 40
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9265 0 0
2
44974.7 29
0
14 Logic Display~
6 815 1032 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
44974.7 30
0
14 Logic Display~
6 817 957 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
44974.7 31
0
14 Logic Display~
6 816 904 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
5.90066e-315 5.34643e-315
0
14 NO PushButton~
191 229 834 0 2 5
0 42 31
0
0 0 4704 0
0
2 S2
-7 -22 7 -14
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9281 0 0
2
5.90066e-315 5.36716e-315
0
5 4049~
219 202 386 0 2 22
0 42 44
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
8464 0 0
2
5.90066e-315 5.37752e-315
0
9 2-In AND~
219 224 427 0 3 22
0 44 35 43
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7168 0 0
2
5.90066e-315 5.38788e-315
0
5 4049~
219 190 297 0 2 22
0 47 46
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3171 0 0
2
5.90066e-315 5.39306e-315
0
7 Ground~
168 357 1484 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4139 0 0
2
5.90066e-315 5.39824e-315
0
2 +V
167 163 761 0 1 3
0 31
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
5.90066e-315 5.40342e-315
0
14 NO PushButton~
191 227 794 0 2 5
0 47 31
0
0 0 4704 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5283 0 0
2
5.90066e-315 5.4086e-315
0
8 3-In OR~
219 299 352 0 4 22
0 45 40 43 48
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
6874 0 0
2
5.90066e-315 5.41378e-315
0
9 2-In AND~
219 220 350 0 3 22
0 46 4 45
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5305 0 0
2
5.90066e-315 5.41896e-315
0
7 Ground~
168 864 600 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
34 0 0
2
5.90066e-315 5.42414e-315
0
4 LED~
171 949 545 0 2 2
10 49 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D13
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
969 0 0
2
5.90066e-315 5.42933e-315
0
4 LED~
171 908 540 0 2 2
10 50 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D12
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8402 0 0
2
5.90066e-315 5.43192e-315
0
4 LED~
171 856 539 0 2 2
10 51 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D11
20 -10 41 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3751 0 0
2
5.90066e-315 5.43451e-315
0
4 LED~
171 802 541 0 2 2
10 37 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D10
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4292 0 0
2
5.90066e-315 5.4371e-315
0
4 LED~
171 744 535 0 2 2
10 41 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D9
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6118 0 0
2
5.90066e-315 5.43969e-315
0
4 LED~
171 685 535 0 2 2
10 35 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
34 0 0
2
5.90066e-315 5.44228e-315
0
4 LED~
171 625 534 0 2 2
10 4 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6357 0 0
2
5.90066e-315 5.44487e-315
0
4 LED~
171 568 532 0 2 2
10 52 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
319 0 0
2
5.90066e-315 5.44746e-315
0
4 LED~
171 509 531 0 2 2
10 53 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3976 0 0
2
5.90066e-315 5.45005e-315
0
4 4017
219 434 448 0 14 29
0 48 36 37 53 52 4 35 41 37
51 50 49 54 94
0
0 0 6880 0
4 4017
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
7634 0 0
2
5.90066e-315 5.45264e-315
0
7 Ground~
168 940 271 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
523 0 0
2
5.90066e-315 5.45523e-315
0
7 Pulser~
4 40 35 0 10 12
0 95 96 5 97 0 0 100 100 6
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6748 0 0
2
5.90066e-315 5.45782e-315
0
9 2-In AND~
219 192 163 0 3 22
0 5 52 56
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6901 0 0
2
44974.7 32
0
4 LED~
171 895 231 0 2 2
10 16 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
842 0 0
2
44974.7 33
0
4 LED~
171 834 229 0 2 2
10 17 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3277 0 0
2
44974.7 34
0
4 LED~
171 776 227 0 2 2
10 18 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4212 0 0
2
44974.7 35
0
4 LED~
171 716 223 0 2 2
10 19 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4720 0 0
2
44974.7 36
0
7 74LS175
131 652 147 0 14 29
0 60 56 59 58 57 55 19 98 18
99 17 100 16 101
0
0 0 4832 0
7 74LS175
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 9 13 12 5 4 15 14 10
11 7 6 2 3 1 9 13 12 5
4 15 14 10 11 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
5551 0 0
2
44974.7 37
0
2 +V
167 503 30 0 1 3
0 60
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6986 0 0
2
44974.7 38
0
7 Ground~
168 268 194 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8745 0 0
2
44974.7 39
0
7 74LS161
96 377 86 0 14 29
0 60 60 5 2 2 2 2 60 60
102 55 57 58 59
0
0 0 6880 0
8 74LS161A
-28 -60 28 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9592 0 0
2
44974.7 40
0
9 Resistor~
219 1410 383 0 3 5
0 25 24 1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8748 0 0
2
44974.7 41
0
9 Resistor~
219 1406 321 0 3 5
0 25 26 1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
44974.7 42
0
9 Resistor~
219 1404 237 0 3 5
0 25 27 1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
631 0 0
2
44974.7 43
0
9 Resistor~
219 1388 156 0 4 5
0 28 25 0 1
0
0 0 864 90
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9466 0 0
2
44974.7 44
0
9 Resistor~
219 275 1140 0 4 5
0 30 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R2
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3266 0 0
2
44974.7 45
0
9 Resistor~
219 282 879 0 4 5
0 38 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R4
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7693 0 0
2
44974.7 46
0
9 Resistor~
219 280 841 0 4 5
0 42 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R3
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3723 0 0
2
5.90066e-315 5.46041e-315
0
9 Resistor~
219 275 803 0 4 5
0 47 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R1
-9 -24 5 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3440 0 0
2
44974.7 47
0
178
2 1 3 0 0 8320 0 1 10 0 0 5
913 799
1275 799
1275 68
1983 68
1983 326
0 1 4 0 0 4096 0 0 1 92 0 3
850 977
850 799
877 799
0 2 5 0 0 4224 0 0 10 93 0 5
1138 924
1138 82
1911 82
1911 335
1989 335
1 0 6 0 0 4224 0 2 0 0 19 2
1903 204
1903 292
1 0 7 0 0 4096 0 3 0 0 18 2
1924 251
1924 283
1 0 8 0 0 4096 0 5 0 0 17 2
1942 255
1942 274
1 0 9 0 0 4096 0 4 0 0 16 2
1960 250
1960 265
13 1 10 0 0 8320 0 10 6 0 0 4
2053 380
2079 380
2079 470
2123 470
11 1 11 0 0 8320 0 10 7 0 0 4
2053 362
2085 362
2085 421
2122 421
9 1 12 0 0 4224 0 10 8 0 0 4
2053 344
2102 344
2102 377
2121 377
7 1 13 0 0 8320 0 10 9 0 0 3
2053 326
2053 332
2109 332
13 0 9 0 0 8192 0 12 0 0 16 4
1906 429
1927 429
1927 342
1978 342
14 0 8 0 0 8192 0 12 0 0 17 3
1906 438
1974 438
1974 361
15 0 7 0 0 4096 0 12 0 0 18 3
1906 447
1985 447
1985 371
16 0 6 0 0 0 0 12 0 0 19 3
1906 456
1980 456
1980 380
3 13 9 0 0 8320 0 10 13 0 0 4
1989 353
1978 353
1978 265
1895 265
14 4 8 0 0 8320 0 13 10 0 0 4
1895 274
1974 274
1974 362
1989 362
15 5 7 0 0 8320 0 13 10 0 0 4
1895 283
1965 283
1965 371
1989 371
16 6 6 0 0 0 0 13 10 0 0 4
1895 292
1959 292
1959 380
1989 380
2 17 14 0 0 4224 0 11 12 0 0 2
1780 384
1836 384
1 0 15 0 0 12288 0 11 0 0 76 4
1744 384
1723 384
1723 405
1795 405
17 0 15 0 0 0 0 13 0 0 76 2
1825 220
1795 220
5 0 16 0 0 4224 0 12 0 0 160 3
1842 429
1062 429
1062 174
6 0 17 0 0 4224 0 12 0 0 161 3
1842 438
1054 438
1054 156
7 0 18 0 0 4224 0 12 0 0 162 3
1842 447
1047 447
1047 138
8 0 19 0 0 4224 0 12 0 0 163 3
1842 456
1040 456
1040 120
5 0 20 0 0 8320 0 13 0 0 35 4
1831 265
1750 265
1750 168
1695 168
6 0 21 0 0 4224 0 13 0 0 31 4
1831 274
1739 274
1739 218
1697 218
7 0 22 0 0 12416 0 13 0 0 34 4
1831 283
1793 283
1793 287
1696 287
8 0 23 0 0 8320 0 13 0 0 33 3
1831 292
1831 327
1697 327
1 11 21 0 0 0 0 16 25 0 0 5
1697 207
1697 218
1682 218
1682 202
1668 202
2 0 24 0 0 8192 0 70 0 0 47 3
1392 383
1387 383
1387 330
1 11 23 0 0 0 0 14 24 0 0 5
1697 323
1697 327
1681 327
1681 321
1667 321
1 9 22 0 0 0 0 15 24 0 0 5
1696 283
1696 287
1681 287
1681 285
1667 285
1 9 20 0 0 0 0 17 25 0 0 5
1695 164
1695 168
1682 168
1682 166
1668 166
1 0 25 0 0 4096 0 70 0 0 64 2
1428 383
1457 383
1 0 25 0 0 4096 0 71 0 0 51 2
1424 321
1458 321
2 0 26 0 0 4096 0 71 0 0 48 2
1388 321
1388 294
1 0 25 0 0 4096 0 72 0 0 64 2
1422 237
1457 237
2 0 27 0 0 4096 0 72 0 0 49 2
1386 237
1386 211
2 0 25 0 0 4096 0 73 0 0 64 2
1388 138
1457 138
1 0 28 0 0 4096 0 73 0 0 50 2
1388 174
1388 175
2 0 2 0 0 12288 0 19 0 0 63 4
1321 330
1268 330
1268 358
1513 358
2 0 2 0 0 0 0 18 0 0 63 4
1320 294
1269 294
1269 257
1513 257
2 0 2 0 0 0 0 20 0 0 63 4
1322 211
1270 211
1270 249
1513 249
2 0 2 0 0 0 0 21 0 0 63 4
1323 175
1272 175
1272 124
1513 124
1 7 24 0 0 4224 0 19 24 0 0 2
1355 330
1597 330
3 1 26 0 0 4224 0 24 18 0 0 2
1597 294
1354 294
7 1 27 0 0 4224 0 25 20 0 0 2
1598 211
1356 211
1 3 28 0 0 4224 0 21 25 0 0 2
1357 175
1598 175
6 0 25 0 0 4096 0 24 0 0 64 2
1603 321
1457 321
5 0 25 0 0 0 0 24 0 0 64 2
1603 312
1457 312
2 0 25 0 0 0 0 24 0 0 64 2
1603 285
1457 285
1 0 25 0 0 0 0 24 0 0 64 2
1603 276
1457 276
6 0 25 0 0 4096 0 25 0 0 64 2
1604 202
1457 202
5 0 25 0 0 0 0 25 0 0 64 2
1604 193
1457 193
2 0 25 0 0 0 0 25 0 0 64 2
1604 166
1457 166
1 0 25 0 0 0 0 25 0 0 64 2
1604 157
1457 157
4 0 25 0 0 0 0 24 0 0 64 2
1597 303
1457 303
4 0 25 0 0 0 0 25 0 0 64 2
1598 184
1457 184
8 0 25 0 0 0 0 24 0 0 64 2
1597 339
1457 339
8 0 25 0 0 0 0 25 0 0 64 2
1598 220
1457 220
1 0 2 0 0 8320 0 22 0 0 0 3
1541 21
1513 21
1513 1729
1 0 25 0 0 4224 0 23 0 0 0 2
1457 55
1457 1729
0 0 2 0 0 0 0 0 0 0 107 4
1227 887
466 887
466 1014
357 1014
2 1 29 0 0 4224 0 26 31 0 0 4
293 1033
494 1033
494 1183
514 1183
0 1 4 0 0 4096 0 0 26 92 0 7
665 841
400 841
400 984
221 984
221 1032
257 1032
257 1033
2 0 30 0 0 12416 0 31 0 0 70 5
520 1192
444 1192
444 1050
245 1050
245 1140
2 0 2 0 0 0 0 74 0 0 107 2
293 1140
357 1140
1 1 30 0 0 0 0 27 74 0 0 3
230 1139
230 1140
257 1140
2 0 31 0 0 4096 0 27 0 0 110 2
196 1139
163 1139
1 0 32 0 0 4096 0 28 0 0 75 2
813 1295
813 1296
1 0 15 0 0 0 0 29 0 0 76 2
812 1208
812 1210
1 0 33 0 0 4096 0 30 0 0 77 2
815 1111
815 1114
4 0 32 0 0 12416 0 31 0 0 0 4
584 1219
676 1219
676 1296
1142 1296
5 0 15 0 0 4224 0 31 0 0 0 3
584 1210
1795 1210
1795 24
6 0 33 0 0 12416 0 31 0 0 0 4
584 1201
677 1201
677 1114
1142 1114
7 3 34 0 0 12416 0 31 31 0 0 6
584 1192
627 1192
627 1082
470 1082
470 1210
520 1210
0 0 35 0 0 4096 0 0 0 136 94 2
721 475
721 915
2 2 36 0 0 4224 0 32 58 0 0 2
299 475
402 475
0 3 37 0 0 8320 0 0 58 138 0 5
824 457
824 619
350 619
350 493
402 493
0 1 38 0 0 12416 0 0 34 85 0 5
256 880
256 851
107 851
107 527
214 527
2 0 31 0 0 4096 0 33 0 0 110 2
212 879
163 879
2 0 2 0 0 0 0 75 0 0 107 4
300 879
353 879
353 881
358 881
1 1 38 0 0 0 0 33 75 0 0 5
246 879
246 880
256 880
256 879
264 879
2 1 39 0 0 12416 0 34 35 0 0 6
250 527
265 527
265 547
208 547
208 558
216 558
3 2 40 0 0 8320 0 35 46 0 0 6
261 567
326 567
326 392
260 392
260 352
287 352
0 2 41 0 0 12288 0 0 35 90 0 6
616 799
481 799
481 625
211 625
211 576
216 576
1 0 41 0 0 0 0 36 0 0 90 2
815 1050
815 1050
0 0 41 0 0 16512 0 0 0 137 0 5
767 466
767 799
611 799
611 1050
1141 1050
1 0 4 0 0 0 0 37 0 0 92 4
817 975
817 976
813 976
813 977
0 0 4 0 0 8192 0 0 0 112 0 3
665 709
665 977
1140 977
0 0 5 0 0 0 0 0 0 0 0 4
816 924
1192 924
1192 914
1227 914
0 0 35 0 0 0 0 0 0 0 0 2
747 915
709 915
0 2 35 0 0 0 0 0 41 79 0 5
721 879
435 879
435 655
200 655
200 436
1 0 42 0 0 8320 0 40 0 0 98 5
187 386
130 386
130 820
255 820
255 841
2 0 2 0 0 0 0 76 0 0 107 2
298 841
358 841
1 1 42 0 0 0 0 39 76 0 0 3
246 842
246 841
262 841
2 0 31 0 0 0 0 39 0 0 110 2
212 842
163 842
3 3 43 0 0 8320 0 41 46 0 0 4
245 427
283 427
283 361
286 361
2 1 44 0 0 12416 0 40 41 0 0 6
223 386
250 386
250 401
193 401
193 418
200 418
1 3 45 0 0 4224 0 46 47 0 0 4
286 343
254 343
254 350
241 350
1 0 5 0 0 0 0 32 0 0 148 2
263 475
91 475
2 1 46 0 0 8320 0 42 47 0 0 5
211 297
211 315
179 315
179 341
196 341
0 1 47 0 0 12416 0 0 42 108 0 5
251 803
251 729
120 729
120 297
175 297
2 0 2 0 0 0 0 77 0 0 107 2
293 803
358 803
1 0 2 0 0 0 0 43 0 0 0 4
357 1478
357 881
358 881
358 749
1 1 47 0 0 0 0 45 77 0 0 3
244 802
244 803
257 803
2 0 31 0 0 0 0 45 0 0 110 2
210 802
163 802
1 0 31 0 0 4224 0 44 0 0 0 2
163 770
163 1469
4 1 48 0 0 8320 0 46 58 0 0 4
332 352
391 352
391 466
396 466
2 0 4 0 0 12416 0 47 0 0 135 5
196 359
177 359
177 709
665 709
665 484
1 0 2 0 0 0 0 48 0 0 132 2
864 594
864 570
2 0 2 0 0 0 0 49 0 0 115 4
949 555
949 560
899 560
899 565
2 0 2 0 0 0 0 50 0 0 132 4
908 550
908 565
887 565
887 570
2 0 2 0 0 0 0 51 0 0 132 2
856 549
856 570
1 0 49 0 0 4096 0 49 0 0 141 4
949 535
949 435
922 435
922 430
1 0 50 0 0 4096 0 50 0 0 140 2
908 530
908 439
1 0 51 0 0 4096 0 51 0 0 139 2
856 529
856 448
1 0 37 0 0 0 0 52 0 0 138 2
802 531
802 457
1 0 41 0 0 0 0 53 0 0 137 2
744 525
744 466
1 0 35 0 0 0 0 54 0 0 136 2
685 525
685 475
1 0 4 0 0 0 0 55 0 0 135 2
625 524
625 484
1 0 52 0 0 4096 0 56 0 0 134 2
568 522
568 493
1 0 53 0 0 4096 0 57 0 0 133 2
509 521
509 502
2 0 2 0 0 0 0 52 0 0 132 2
802 551
802 570
2 0 2 0 0 0 0 53 0 0 132 2
744 545
744 570
2 0 2 0 0 0 0 54 0 0 132 2
685 545
685 570
2 0 2 0 0 0 0 55 0 0 132 2
625 544
625 570
2 0 2 0 0 0 0 56 0 0 132 2
568 542
568 570
2 0 2 0 0 0 0 57 0 0 132 2
509 541
509 570
0 0 2 0 0 0 0 0 0 0 0 2
482 570
894 570
4 0 53 0 0 4224 0 58 0 0 0 2
466 502
946 502
5 0 52 0 0 4096 0 58 0 0 0 2
466 493
959 493
6 0 4 0 0 0 0 58 0 0 0 2
466 484
947 484
7 0 35 0 0 4224 0 58 0 0 0 2
466 475
940 475
8 0 41 0 0 0 0 58 0 0 0 2
466 466
945 466
9 0 37 0 0 0 0 58 0 0 0 2
466 457
935 457
10 0 51 0 0 4224 0 58 0 0 0 2
466 448
940 448
11 0 50 0 0 4224 0 58 0 0 0 2
466 439
934 439
12 0 49 0 0 4224 0 58 0 0 0 2
466 430
929 430
13 0 54 0 0 4224 0 58 0 0 0 3
466 421
926 421
926 424
2 0 2 0 0 0 0 62 0 0 147 2
895 241
895 265
2 0 2 0 0 0 0 63 0 0 147 2
834 239
834 265
2 0 2 0 0 0 0 64 0 0 147 2
776 237
776 265
2 0 2 0 0 0 0 65 0 0 147 2
716 233
716 265
1 0 2 0 0 0 0 59 0 0 0 2
940 265
692 265
0 0 5 0 0 0 0 0 0 150 0 2
91 457
91 987
3 0 5 0 0 0 0 69 0 0 150 2
345 68
91 68
3 0 5 0 0 0 0 60 0 0 0 4
64 26
91 26
91 459
107 459
6 0 55 0 0 4096 0 66 0 0 152 2
620 174
527 174
11 0 55 0 0 4224 0 69 0 0 0 3
409 95
527 95
527 199
2 0 52 0 0 16512 0 61 0 0 134 7
168 172
158 172
158 171
150 171
150 680
587 680
587 493
1 0 5 0 0 0 0 61 0 0 150 5
168 154
168 127
237 127
237 80
91 80
2 3 56 0 0 12416 0 66 61 0 0 6
620 129
555 129
555 258
235 258
235 163
213 163
1 0 16 0 0 0 0 62 0 0 160 2
895 221
895 174
1 0 17 0 0 0 0 63 0 0 161 2
834 219
834 156
1 0 18 0 0 0 0 64 0 0 162 2
776 217
776 138
1 0 19 0 0 0 0 65 0 0 163 2
716 213
716 120
13 0 16 0 0 0 0 66 0 0 0 2
684 174
1226 174
11 0 17 0 0 0 0 66 0 0 0 2
684 156
1223 156
9 0 18 0 0 0 0 66 0 0 0 2
684 138
1224 138
7 0 19 0 0 0 0 66 0 0 0 2
684 120
1225 120
5 0 57 0 0 4224 0 66 0 0 172 2
620 165
479 165
4 0 58 0 0 4224 0 66 0 0 173 2
620 156
413 156
3 0 59 0 0 4224 0 66 0 0 174 2
620 147
355 147
1 0 60 0 0 12288 0 66 0 0 171 6
614 120
597 120
597 55
507 55
507 50
495 50
1 0 60 0 0 0 0 69 0 0 169 3
345 50
330 50
330 7
2 0 60 0 0 12416 0 69 0 0 171 5
345 59
309 59
309 7
461 7
461 50
9 0 60 0 0 0 0 69 0 0 171 3
415 59
489 59
489 50
8 1 60 0 0 0 0 69 67 0 0 4
415 50
495 50
495 39
503 39
0 12 57 0 0 0 0 0 69 0 0 3
479 172
479 104
409 104
0 13 58 0 0 0 0 0 69 0 0 5
413 172
413 141
428 141
428 113
409 113
0 14 59 0 0 0 0 0 69 0 0 5
355 169
355 136
423 136
423 122
409 122
0 1 2 0 0 0 0 0 68 176 0 5
345 118
262 118
262 175
268 175
268 188
7 6 2 0 0 0 0 69 69 0 0 2
345 122
345 113
5 6 2 0 0 0 0 69 69 0 0 2
345 104
345 113
4 5 2 0 0 0 0 69 69 0 0 2
345 95
345 104
15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
1577 38 1746 53
1591 50 1731 61
20 Venn Diagram Circuit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
435 818 649 841
447 828 636 843
27 Question Mode Change Enable
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 38
1155 1275 1448 1298
1168 1285 1434 1300
38 To master/slave selector of Expression
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
1148 1191 1455 1214
1161 1201 1441 1216
40 To master/slave selector of Venn Diagram
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
901 1269 1061 1292
914 1279 1047 1294
19 Expression Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
900 1182 1073 1205
912 1192 1060 1207
21 Venn Diagram Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
901 1084 984 1107
914 1094 970 1109
8 DIY Mode
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
477 655 630 678
490 665 616 680
18 Load Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
-11 68 100 91
2 78 86 93
12 Clock Signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
459 327 605 350
472 337 591 352
17 Master Controller
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
870 1016 1035 1039
882 1026 1022 1041
20 Output Enable signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
871 86 987 109
883 96 974 111
13 Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
610 10 796 33
622 20 783 35
23 Random Number Generator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
871 948 1050 971
883 958 1037 973
22 Reset signal for slave
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
870 893 1049 916
882 903 1036 918
22 Master Clock for Slave
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
