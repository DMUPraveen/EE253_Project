CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 250 30 90 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 D:\Programs\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.209790 0.500000
855 80 1534 795
9437202 0
0
6 Title:
5 Name:
0
0
0
58
13 Logic Switch~
5 1170 1098 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -19 8 -11
2 V7
-6 -24 8 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
523 0 0
2
44971.5 0
0
13 Logic Switch~
5 1170 1064 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -18 8 -10
2 V6
-6 -24 8 -16
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6748 0 0
2
44971.5 0
0
13 Logic Switch~
5 1169 1032 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6901 0 0
2
44971.5 0
0
13 Logic Switch~
5 1168 999 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -17 8 -9
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
842 0 0
2
44971.5 0
0
14 Logic Display~
6 1375 1085 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
44971.5 0
0
14 Logic Display~
6 1372 1025 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
44971.5 0
0
14 Logic Display~
6 1367 958 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
44971.5 0
0
14 Logic Display~
6 1362 908 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
44971.5 0
0
7 74LS173
129 1259 914 0 14 29
0 2 2 2 27 10 9 8 7 2
2 6 5 4 3
0
0 0 13040 0
7 74LS173
-24 -51 25 -43
2 U9
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 18
65 0 0 0 1 0 0 0
1 U
6986 0 0
2
44971.5 0
0
5 4049~
219 272 1033 0 2 22
0 13 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
8745 0 0
2
44971.5 0
0
14 NO PushButton~
191 213 1131 0 2 5
0 14 15
0
0 0 4720 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9592 0 0
2
44971.5 0
0
14 Logic Display~
6 813 1277 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
44971.5 0
0
14 Logic Display~
6 812 1190 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
44971.5 0
0
14 Logic Display~
6 815 1093 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
44971.5 0
0
4 4017
219 552 1165 0 14 29
0 11 14 19 16 17 18 19 52 53
54 55 56 57 58
0
0 0 6896 0
4 4017
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
9466 0 0
2
44971.4 0
0
5 4049~
219 278 475 0 2 22
0 28 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
3266 0 0
2
44971.4 0
0
14 NO PushButton~
191 229 871 0 2 5
0 23 15
0
0 0 4720 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7693 0 0
2
44971.4 0
0
5 4049~
219 229 527 0 2 22
0 23 24
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
3723 0 0
2
44971.4 0
0
9 2-In AND~
219 240 567 0 3 22
0 24 26 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3440 0 0
2
44971.4 0
0
14 Logic Display~
6 815 1032 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6263 0 0
2
44971.4 0
0
14 Logic Display~
6 817 957 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4900 0 0
2
44971.4 0
0
14 Logic Display~
6 816 904 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8783 0 0
2
5.90066e-315 0
0
9 2-In AND~
219 771 924 0 3 22
0 20 28 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3221 0 0
2
5.90066e-315 0
0
14 NO PushButton~
191 229 834 0 2 5
0 29 15
0
0 0 4720 0
0
2 S2
-7 -22 7 -14
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3215 0 0
2
5.90066e-315 0
0
5 4049~
219 202 386 0 2 22
0 29 31
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
7903 0 0
2
5.90066e-315 0
0
9 2-In AND~
219 224 427 0 3 22
0 31 20 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7121 0 0
2
5.90066e-315 0
0
5 4049~
219 190 297 0 2 22
0 34 33
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
4484 0 0
2
5.90066e-315 0
0
7 Ground~
168 357 1484 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5996 0 0
2
5.90066e-315 0
0
2 +V
167 163 761 0 1 3
0 15
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7804 0 0
2
5.90066e-315 0
0
14 NO PushButton~
191 227 794 0 2 5
0 34 15
0
0 0 4720 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5523 0 0
2
5.90066e-315 0
0
8 3-In OR~
219 299 352 0 4 22
0 32 25 30 35
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3330 0 0
2
5.90066e-315 0
0
9 2-In AND~
219 220 350 0 3 22
0 33 13 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3465 0 0
2
5.90066e-315 0
0
7 Ground~
168 864 600 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8396 0 0
2
5.90066e-315 0
0
4 LED~
171 949 545 0 2 2
10 36 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D13
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3685 0 0
2
5.90066e-315 0
0
4 LED~
171 908 540 0 2 2
10 37 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D12
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7849 0 0
2
5.90066e-315 0
0
4 LED~
171 856 539 0 2 2
10 38 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D11
20 -10 41 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6343 0 0
2
5.90066e-315 0
0
4 LED~
171 802 541 0 2 2
10 22 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D10
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7376 0 0
2
5.90066e-315 0
0
4 LED~
171 744 535 0 2 2
10 26 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D9
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9156 0 0
2
5.90066e-315 0
0
4 LED~
171 685 535 0 2 2
10 20 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5776 0 0
2
5.90066e-315 0
0
4 LED~
171 625 534 0 2 2
10 13 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7207 0 0
2
5.90066e-315 0
0
4 LED~
171 568 532 0 2 2
10 39 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4459 0 0
2
5.90066e-315 0
0
4 LED~
171 509 531 0 2 2
10 40 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3760 0 0
2
5.90066e-315 0
0
4 4017
219 434 448 0 14 29
0 35 21 22 40 39 13 20 26 22
38 37 36 41 59
0
0 0 6896 0
4 4017
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
754 0 0
2
5.90066e-315 0
0
7 Ground~
168 940 271 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9767 0 0
2
5.90066e-315 0
0
7 Pulser~
4 40 35 0 10 12
0 60 61 28 62 0 0 5 5 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7978 0 0
2
5.90066e-315 0
0
9 2-In AND~
219 192 163 0 3 22
0 28 39 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3142 0 0
2
44971.4 0
0
4 LED~
171 895 231 0 2 2
10 44 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3284 0 0
2
44971.4 1
0
4 LED~
171 834 229 0 2 2
10 45 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
659 0 0
2
44971.4 2
0
4 LED~
171 776 227 0 2 2
10 46 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3800 0 0
2
44971.4 3
0
4 LED~
171 716 223 0 2 2
10 47 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6792 0 0
2
44971.4 4
0
7 74LS175
131 652 147 0 14 29
0 51 43 50 49 48 42 47 63 46
64 45 65 44 66
0
0 0 4848 0
7 74LS175
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 9 13 12 5 4 15 14 10
11 7 6 2 3 1 9 13 12 5
4 15 14 10 11 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3701 0 0
2
44971.4 5
0
2 +V
167 503 30 0 1 3
0 51
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6316 0 0
2
44971.4 6
0
7 Ground~
168 268 194 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8734 0 0
2
44971.4 7
0
7 74LS161
96 377 86 0 14 29
0 51 51 28 2 2 2 2 51 51
67 42 48 49 50
0
0 0 6896 0
8 74LS161A
-28 -60 28 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
7988 0 0
2
44971.4 8
0
9 Resistor~
219 275 1140 0 4 5
0 14 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3217 0 0
2
44971.5 0
0
9 Resistor~
219 282 879 0 4 5
0 23 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R4
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3965 0 0
2
44971.4 0
0
9 Resistor~
219 280 841 0 4 5
0 29 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8239 0 0
2
5.90066e-315 0
0
9 Resistor~
219 275 803 0 4 5
0 34 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-9 -24 5 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
828 0 0
2
44971.4 9
0
128
14 1 3 0 0 8320 0 9 5 0 0 4
1291 950
1303 950
1303 1103
1375 1103
13 1 4 0 0 8320 0 9 6 0 0 4
1291 941
1313 941
1313 1043
1372 1043
12 1 5 0 0 8320 0 9 7 0 0 4
1291 932
1326 932
1326 976
1367 976
1 11 6 0 0 4224 0 8 9 0 0 5
1362 926
1309 926
1309 914
1291 914
1291 923
1 8 7 0 0 8320 0 1 9 0 0 3
1182 1098
1227 1098
1227 950
7 1 8 0 0 8320 0 9 2 0 0 4
1227 941
1219 941
1219 1064
1182 1064
1 6 9 0 0 8320 0 3 9 0 0 4
1181 1032
1214 1032
1214 932
1227 932
1 5 10 0 0 8320 0 4 9 0 0 4
1180 999
1203 999
1203 923
1227 923
9 0 2 0 0 8192 0 9 0 0 12 4
1297 887
1297 850
1138 850
1138 887
9 10 2 0 0 0 0 9 9 0 0 2
1297 887
1297 896
2 0 2 0 0 0 0 9 0 0 12 3
1221 896
1187 896
1187 887
1 0 2 0 0 4224 0 9 0 0 57 4
1227 887
466 887
466 1014
357 1014
3 2 2 0 0 0 0 9 9 0 0 2
1221 905
1221 896
2 1 11 0 0 4224 0 10 15 0 0 4
293 1033
494 1033
494 1183
514 1183
0 1 13 0 0 4096 0 0 10 40 0 7
665 841
400 841
400 984
221 984
221 1032
257 1032
257 1033
2 0 14 0 0 12416 0 15 0 0 18 5
520 1192
444 1192
444 1050
245 1050
245 1140
2 0 2 0 0 0 0 55 0 0 57 2
293 1140
357 1140
1 1 14 0 0 0 0 11 55 0 0 3
230 1139
230 1140
257 1140
2 0 15 0 0 4096 0 11 0 0 60 2
196 1139
163 1139
1 0 16 0 0 4096 0 12 0 0 23 2
813 1295
813 1296
1 0 17 0 0 4096 0 13 0 0 24 2
812 1208
812 1210
1 0 18 0 0 4096 0 14 0 0 25 2
815 1111
815 1114
4 0 16 0 0 12416 0 15 0 0 0 4
584 1219
676 1219
676 1296
1142 1296
5 0 17 0 0 4224 0 15 0 0 0 2
584 1210
1144 1210
6 0 18 0 0 12416 0 15 0 0 0 4
584 1201
677 1201
677 1114
1142 1114
7 3 19 0 0 12416 0 15 15 0 0 6
584 1192
627 1192
627 1082
470 1082
470 1210
520 1210
0 0 20 0 0 4096 0 0 0 86 44 2
721 475
721 915
2 2 21 0 0 4224 0 16 43 0 0 2
299 475
402 475
0 3 22 0 0 8320 0 0 43 88 0 5
824 457
824 619
350 619
350 493
402 493
0 1 23 0 0 12416 0 0 18 33 0 5
256 880
256 851
107 851
107 527
214 527
2 0 15 0 0 4096 0 17 0 0 60 2
212 879
163 879
2 0 2 0 0 0 0 56 0 0 57 4
300 879
353 879
353 881
358 881
1 1 23 0 0 0 0 17 56 0 0 5
246 879
246 880
256 880
256 879
264 879
2 1 24 0 0 12416 0 18 19 0 0 6
250 527
265 527
265 547
208 547
208 558
216 558
3 2 25 0 0 8320 0 19 31 0 0 6
261 567
326 567
326 392
260 392
260 352
287 352
0 2 26 0 0 12288 0 0 19 38 0 6
616 799
481 799
481 625
211 625
211 576
216 576
1 0 26 0 0 0 0 20 0 0 38 2
815 1050
815 1050
0 0 26 0 0 16512 0 0 0 87 0 5
767 466
767 799
611 799
611 1050
1141 1050
1 0 13 0 0 0 0 21 0 0 40 4
817 975
817 976
813 976
813 977
0 0 13 0 0 8192 0 0 0 62 0 3
665 709
665 977
1140 977
0 4 27 0 0 4224 0 0 9 42 0 4
816 924
1192 924
1192 914
1227 914
1 3 27 0 0 128 0 22 23 0 0 3
816 922
816 924
792 924
2 0 28 0 0 4224 0 23 0 0 98 2
747 933
91 933
1 0 20 0 0 0 0 23 0 0 0 2
747 915
709 915
0 2 20 0 0 128 0 0 26 27 0 5
721 879
435 879
435 655
200 655
200 436
1 0 29 0 0 8320 0 25 0 0 48 5
187 386
130 386
130 820
255 820
255 841
2 0 2 0 0 0 0 57 0 0 57 2
298 841
358 841
1 1 29 0 0 0 0 24 57 0 0 3
246 842
246 841
262 841
2 0 15 0 0 0 0 24 0 0 60 2
212 842
163 842
3 3 30 0 0 8320 0 26 31 0 0 4
245 427
283 427
283 361
286 361
2 1 31 0 0 12416 0 25 26 0 0 6
223 386
250 386
250 401
193 401
193 418
200 418
1 3 32 0 0 4224 0 31 32 0 0 4
286 343
254 343
254 350
241 350
1 0 28 0 0 0 0 16 0 0 98 2
263 475
91 475
2 1 33 0 0 8320 0 27 32 0 0 5
211 297
211 315
179 315
179 341
196 341
0 1 34 0 0 12416 0 0 27 58 0 5
251 803
251 729
120 729
120 297
175 297
2 0 2 0 0 0 0 58 0 0 57 2
293 803
358 803
1 0 2 0 0 128 0 28 0 0 0 4
357 1478
357 881
358 881
358 749
1 1 34 0 0 0 0 30 58 0 0 3
244 802
244 803
257 803
2 0 15 0 0 0 0 30 0 0 60 2
210 802
163 802
1 0 15 0 0 4224 0 29 0 0 0 2
163 770
163 1469
4 1 35 0 0 8320 0 31 43 0 0 4
332 352
391 352
391 466
396 466
2 0 13 0 0 12416 0 32 0 0 85 5
196 359
177 359
177 709
665 709
665 484
1 0 2 0 0 0 0 33 0 0 82 2
864 594
864 570
2 0 2 0 0 0 0 34 0 0 65 4
949 555
949 560
899 560
899 565
2 0 2 0 0 0 0 35 0 0 82 4
908 550
908 565
887 565
887 570
2 0 2 0 0 0 0 36 0 0 82 2
856 549
856 570
1 0 36 0 0 4096 0 34 0 0 91 4
949 535
949 435
922 435
922 430
1 0 37 0 0 4096 0 35 0 0 90 2
908 530
908 439
1 0 38 0 0 4096 0 36 0 0 89 2
856 529
856 448
1 0 22 0 0 0 0 37 0 0 88 2
802 531
802 457
1 0 26 0 0 0 0 38 0 0 87 2
744 525
744 466
1 0 20 0 0 0 0 39 0 0 86 2
685 525
685 475
1 0 13 0 0 0 0 40 0 0 85 2
625 524
625 484
1 0 39 0 0 4096 0 41 0 0 84 2
568 522
568 493
1 0 40 0 0 4096 0 42 0 0 83 2
509 521
509 502
2 0 2 0 0 0 0 37 0 0 82 2
802 551
802 570
2 0 2 0 0 0 0 38 0 0 82 2
744 545
744 570
2 0 2 0 0 0 0 39 0 0 82 2
685 545
685 570
2 0 2 0 0 0 0 40 0 0 82 2
625 544
625 570
2 0 2 0 0 0 0 41 0 0 82 2
568 542
568 570
2 0 2 0 0 0 0 42 0 0 82 2
509 541
509 570
0 0 2 0 0 128 0 0 0 0 0 2
482 570
894 570
4 0 40 0 0 4224 0 43 0 0 0 2
466 502
946 502
5 0 39 0 0 4096 0 43 0 0 0 2
466 493
959 493
6 0 13 0 0 0 0 43 0 0 0 2
466 484
947 484
7 0 20 0 0 4224 0 43 0 0 0 2
466 475
940 475
8 0 26 0 0 128 0 43 0 0 0 2
466 466
945 466
9 0 22 0 0 128 0 43 0 0 0 2
466 457
935 457
10 0 38 0 0 4224 0 43 0 0 0 2
466 448
940 448
11 0 37 0 0 4224 0 43 0 0 0 2
466 439
934 439
12 0 36 0 0 4224 0 43 0 0 0 2
466 430
929 430
13 0 41 0 0 4224 0 43 0 0 0 3
466 421
926 421
926 424
2 0 2 0 0 0 0 47 0 0 97 2
895 241
895 265
2 0 2 0 0 0 0 48 0 0 97 2
834 239
834 265
2 0 2 0 0 0 0 49 0 0 97 2
776 237
776 265
2 0 2 0 0 0 0 50 0 0 97 2
716 233
716 265
1 0 2 0 0 0 0 44 0 0 0 2
940 265
692 265
0 0 28 0 0 0 0 0 0 100 0 2
91 457
91 987
3 0 28 0 0 0 0 54 0 0 100 2
345 68
91 68
3 0 28 0 0 0 0 45 0 0 0 4
64 26
91 26
91 459
107 459
6 0 42 0 0 4096 0 51 0 0 102 2
620 174
527 174
11 0 42 0 0 4224 0 54 0 0 0 3
409 95
527 95
527 199
2 0 39 0 0 16512 0 46 0 0 84 7
168 172
158 172
158 171
150 171
150 680
587 680
587 493
1 0 28 0 0 0 0 46 0 0 100 5
168 154
168 127
237 127
237 80
91 80
2 3 43 0 0 12416 0 51 46 0 0 6
620 129
555 129
555 258
235 258
235 163
213 163
1 0 44 0 0 4096 0 47 0 0 110 2
895 221
895 174
1 0 45 0 0 4096 0 48 0 0 111 2
834 219
834 156
1 0 46 0 0 4096 0 49 0 0 112 2
776 217
776 138
1 0 47 0 0 4096 0 50 0 0 113 2
716 213
716 120
13 0 44 0 0 4224 0 51 0 0 0 2
684 174
999 174
11 0 45 0 0 4224 0 51 0 0 0 2
684 156
989 156
9 0 46 0 0 4224 0 51 0 0 0 2
684 138
975 138
7 0 47 0 0 4224 0 51 0 0 0 2
684 120
961 120
5 0 48 0 0 4224 0 51 0 0 122 2
620 165
479 165
4 0 49 0 0 4224 0 51 0 0 123 2
620 156
413 156
3 0 50 0 0 4224 0 51 0 0 124 2
620 147
355 147
1 0 51 0 0 12288 0 51 0 0 121 6
614 120
597 120
597 55
507 55
507 50
495 50
1 0 51 0 0 0 0 54 0 0 119 3
345 50
330 50
330 7
2 0 51 0 0 12416 0 54 0 0 121 5
345 59
309 59
309 7
461 7
461 50
9 0 51 0 0 0 0 54 0 0 121 3
415 59
489 59
489 50
8 1 51 0 0 0 0 54 52 0 0 4
415 50
495 50
495 39
503 39
0 12 48 0 0 0 0 0 54 0 0 3
479 172
479 104
409 104
0 13 49 0 0 0 0 0 54 0 0 5
413 172
413 141
428 141
428 113
409 113
0 14 50 0 0 0 0 0 54 0 0 5
355 169
355 136
423 136
423 122
409 122
0 1 2 0 0 0 0 0 53 126 0 5
345 118
262 118
262 175
268 175
268 188
7 6 2 0 0 0 0 54 54 0 0 2
345 122
345 113
5 6 2 0 0 0 0 54 54 0 0 2
345 104
345 113
4 5 2 0 0 0 0 54 54 0 0 2
345 95
345 104
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
435 818 649 841
447 828 636 843
27 Question Mode Change Enable
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 38
1155 1275 1448 1298
1168 1285 1434 1300
38 To master/slave selector of Expression
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
1148 1191 1455 1214
1161 1201 1441 1216
40 To master/slave selector of Venn Diagram
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
901 1269 1061 1292
914 1279 1047 1294
19 Expression Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
900 1182 1073 1205
912 1192 1060 1207
21 Venn Diagram Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
901 1084 984 1107
914 1094 970 1109
8 DIY Mode
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
477 655 630 678
490 665 616 680
18 Load Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
-11 68 100 91
2 78 86 93
12 Clock Signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
457 327 603 350
470 337 589 352
17 Master Controller
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
870 1016 1035 1039
882 1026 1022 1041
20 Output Enable signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
871 86 987 109
883 96 974 111
13 Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
610 10 796 33
622 20 783 35
23 Random Number Generator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
871 948 1050 971
883 958 1037 973
22 Reset signal for slave
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
870 893 1049 916
882 903 1036 918
22 Master Clock for Slave
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
