CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 D:\Programs\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.209790 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
211
14 Logic Display~
6 2254 1306 0 1 2
12 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5130 0 0
2
44974.9 0
0
14 Logic Display~
6 2210 1305 0 1 2
12 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
44974.9 1
0
14 Logic Display~
6 2168 1305 0 1 2
12 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
44974.9 2
0
14 Logic Display~
6 2124 1304 0 1 2
12 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
44974.9 3
0
14 Logic Display~
6 2045 1305 0 1 2
15 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N0
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
44974.9 4
0
14 Logic Display~
6 2005 1305 0 1 2
15 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44974.9 5
0
14 Logic Display~
6 1961 1304 0 1 2
15 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
44974.9 6
0
14 Logic Display~
6 1920 1304 0 1 2
15 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
44974.9 7
0
6 74136~
219 2307 1418 0 3 22
0 10 5 21
0
0 0 96 0
7 74LS136
-24 -24 25 -16
3 A2D
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
4747 0 0
2
44974.9 8
0
6 74136~
219 2306 1480 0 3 22
0 9 6 20
0
0 0 96 0
7 74LS136
-24 -24 25 -16
3 A2C
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
972 0 0
2
44974.9 9
0
6 74136~
219 2306 1544 0 3 22
0 8 4 19
0
0 0 96 0
7 74LS136
-24 -24 25 -16
3 A2B
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 19 0
1 U
3472 0 0
2
44974.9 10
0
6 74136~
219 2309 1609 0 3 22
0 7 3 18
0
0 0 96 0
7 74LS136
-24 -24 25 -16
3 A2A
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
9998 0 0
2
44974.9 11
0
8 2-In OR~
219 2402 1451 0 3 22
0 21 20 17
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 A1A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
3536 0 0
2
44974.9 12
0
8 2-In OR~
219 2397 1567 0 3 22
0 19 18 16
0
0 0 96 0
6 74LS32
-21 -24 21 -16
4 U31D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
4597 0 0
2
44974.9 13
0
8 2-In OR~
219 2482 1509 0 3 22
0 17 16 15
0
0 0 96 0
6 74LS32
-21 -24 21 -16
4 U31C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
3835 0 0
2
44974.9 14
0
9 Inverter~
13 2595 1451 0 2 22
0 15 14
0
0 0 96 0
6 74LS04
-21 -19 21 -11
4 U32F
-14 -29 14 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 17 0
1 U
3670 0 0
2
44974.9 15
0
9 2-In AND~
219 2676 1403 0 3 22
0 13 14 12
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 U26D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
5616 0 0
2
44974.9 16
0
9 2-In AND~
219 2677 1572 0 3 22
0 13 15 11
0
0 0 96 0
6 74LS08
-21 -24 21 -16
4 U26C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
9323 0 0
2
44974.9 17
0
14 Logic Display~
6 2669 1268 0 1 2
22 13
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 R27
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
44974.9 18
0
14 Logic Display~
6 2764 1398 0 1 2
10 12
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 R26
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44974.9 19
0
14 Logic Display~
6 2759 1568 0 1 2
14 11
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 R25
14 -26 35 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
44974.9 20
0
8 2-In OR~
219 1094 2430 0 3 22
0 23 22 24
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U31B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
9672 0 0
2
5.90066e-315 0
0
9 Inverter~
13 845 2372 0 2 22
0 46 23
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U32E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 17 0
1 U
7876 0 0
2
5.90066e-315 5.26354e-315
0
9 2-In AND~
219 1224 2804 0 3 22
0 24 48 47
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U26B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
6369 0 0
2
5.90066e-315 5.30499e-315
0
7 Ground~
168 824 2297 0 1 3
0 2
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
5.90066e-315 5.32571e-315
0
9 Inverter~
13 1095 2132 0 2 22
0 62 54
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U32D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 17 0
1 U
7100 0 0
2
5.90066e-315 5.34643e-315
0
9 Inverter~
13 1030 2133 0 2 22
0 63 55
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U32C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 17 0
1 U
3820 0 0
2
5.90066e-315 5.3568e-315
0
9 Inverter~
13 950 2133 0 2 22
0 64 56
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U32B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 17 0
1 U
7678 0 0
2
5.90066e-315 5.36716e-315
0
9 Inverter~
13 887 2132 0 2 22
0 65 57
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U32A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 17 0
1 U
961 0 0
2
5.90066e-315 5.37752e-315
0
9 Inverter~
13 805 2132 0 2 22
0 66 58
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U29F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 14 0
1 U
3178 0 0
2
5.90066e-315 5.38788e-315
0
9 Inverter~
13 744 2133 0 2 22
0 67 59
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U29E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 14 0
1 U
3409 0 0
2
5.90066e-315 5.39306e-315
0
9 Inverter~
13 660 2131 0 2 22
0 68 60
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U29D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 14 0
1 U
3951 0 0
2
5.90066e-315 5.39824e-315
0
9 Inverter~
13 603 2132 0 2 22
0 69 61
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U29C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 14 0
1 U
8885 0 0
2
5.90066e-315 5.40342e-315
0
8 2-In OR~
219 1095 2045 0 3 22
0 27 37 62
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U31A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
3780 0 0
2
5.90066e-315 5.4086e-315
0
8 2-In OR~
219 1030 2042 0 3 22
0 28 38 63
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U30D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
9265 0 0
2
5.90066e-315 5.41378e-315
0
8 2-In OR~
219 946 2041 0 3 22
0 29 39 64
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U30C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
9442 0 0
2
5.90066e-315 5.41896e-315
0
8 2-In OR~
219 889 2041 0 3 22
0 30 40 65
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U30B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
9424 0 0
2
5.90066e-315 5.42414e-315
0
8 2-In OR~
219 806 2043 0 3 22
0 32 42 66
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U30A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
9968 0 0
2
5.90066e-315 5.42933e-315
0
8 2-In OR~
219 743 2045 0 3 22
0 33 43 67
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U18D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
9281 0 0
2
5.90066e-315 5.43192e-315
0
8 2-In OR~
219 662 2045 0 3 22
0 34 44 68
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U18C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
8464 0 0
2
5.90066e-315 5.43451e-315
0
8 2-In OR~
219 600 2047 0 3 22
0 35 45 69
0
0 0 96 270
6 74LS32
-21 -24 21 -16
4 U18B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
7168 0 0
2
5.90066e-315 5.4371e-315
0
7 Ground~
168 623 2332 0 1 3
0 2
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3171 0 0
2
5.90066e-315 5.43969e-315
0
9 Inverter~
13 2376 2641 0 2 22
0 73 89
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U29B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 14 0
1 U
4139 0 0
2
5.90066e-315 5.44228e-315
0
9 Inverter~
13 2411 2637 0 2 22
0 72 88
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U29A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 14 0
1 U
6435 0 0
2
5.90066e-315 5.44487e-315
0
9 Inverter~
13 2443 2638 0 2 22
0 71 87
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U28F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 13 0
1 U
5283 0 0
2
5.90066e-315 5.44746e-315
0
9 Inverter~
13 2476 2637 0 2 22
0 70 86
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U28E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 13 0
1 U
6874 0 0
2
5.90066e-315 5.45005e-315
0
9 Inverter~
13 2207 2641 0 2 22
0 77 93
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U28D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 13 0
1 U
5305 0 0
2
5.90066e-315 5.45264e-315
0
9 Inverter~
13 2242 2637 0 2 22
0 76 92
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U28C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 13 0
1 U
34 0 0
2
5.90066e-315 5.45523e-315
0
9 Inverter~
13 2274 2638 0 2 22
0 75 91
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U28B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 13 0
1 U
969 0 0
2
5.90066e-315 5.45782e-315
0
9 Inverter~
13 2307 2637 0 2 22
0 74 90
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U28A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 13 0
1 U
8402 0 0
2
5.90066e-315 5.46041e-315
0
9 Inverter~
13 2038 2642 0 2 22
0 81 97
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U27F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
3751 0 0
2
5.90066e-315 5.463e-315
0
9 Inverter~
13 2073 2638 0 2 22
0 80 96
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U27E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
4292 0 0
2
5.90066e-315 5.46559e-315
0
9 Inverter~
13 2105 2639 0 2 22
0 79 95
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U27D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
6118 0 0
2
5.90066e-315 5.46818e-315
0
9 Inverter~
13 2138 2638 0 2 22
0 78 94
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U27C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
34 0 0
2
5.90066e-315 5.47077e-315
0
9 Inverter~
13 1974 2642 0 2 22
0 82 98
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U27B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
6357 0 0
2
5.90066e-315 5.47207e-315
0
9 Inverter~
13 1941 2643 0 2 22
0 83 99
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U27A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
319 0 0
2
5.90066e-315 5.47336e-315
0
9 Inverter~
13 1909 2642 0 2 22
0 84 100
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U16F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 5 0
1 U
3976 0 0
2
5.90066e-315 5.47466e-315
0
14 Logic Display~
6 1877 2595 0 1 2
22 101
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L26
-9 -19 12 -11
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
5.90066e-315 5.47595e-315
0
14 Logic Display~
6 1912 2594 0 1 2
10 100
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L25
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
5.90066e-315 5.47725e-315
0
14 Logic Display~
6 1944 2594 0 1 2
10 99
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L24
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
5.90066e-315 5.47854e-315
0
14 Logic Display~
6 1977 2595 0 1 2
10 98
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L23
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
5.90066e-315 5.47984e-315
0
14 Logic Display~
6 2141 2593 0 1 2
10 94
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L22
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
5.90066e-315 5.48113e-315
0
14 Logic Display~
6 2076 2592 0 1 2
10 96
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L21
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
5.90066e-315 5.48243e-315
0
14 Logic Display~
6 2041 2593 0 1 2
10 97
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
5.90066e-315 5.48372e-315
0
14 Logic Display~
6 2309 2592 0 1 2
10 90
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.90066e-315 5.48502e-315
0
14 Logic Display~
6 2276 2591 0 1 2
10 91
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
5.90066e-315 5.48631e-315
0
14 Logic Display~
6 2244 2591 0 1 2
10 92
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
5.90066e-315 5.48761e-315
0
14 Logic Display~
6 2209 2592 0 1 2
10 93
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
5.90066e-315 5.4889e-315
0
14 Logic Display~
6 2478 2592 0 1 2
10 86
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
5.90066e-315 5.4902e-315
0
14 Logic Display~
6 2445 2591 0 1 2
10 87
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.90066e-315 5.49149e-315
0
14 Logic Display~
6 2413 2591 0 1 2
10 88
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90066e-315 5.49279e-315
0
14 Logic Display~
6 2378 2592 0 1 2
10 89
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
5.90066e-315 5.49408e-315
0
14 Logic Display~
6 2108 2592 0 1 2
10 95
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9466 0 0
2
5.90066e-315 5.49538e-315
0
9 Inverter~
13 1874 2646 0 2 22
0 85 101
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U16E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 5 0
1 U
3266 0 0
2
5.90066e-315 5.49667e-315
0
9 Inverter~
13 519 3138 0 2 22
0 22 106
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U16D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
7693 0 0
2
5.90066e-315 5.49797e-315
0
9 2-In AND~
219 991 3060 0 3 22
0 50 25 112
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U26A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3723 0 0
2
5.90066e-315 5.49926e-315
0
8 3-In OR~
219 1087 3049 0 4 22
0 113 112 111 107
0
0 0 608 0
4 4075
-14 -24 14 -16
4 U25B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
3440 0 0
2
5.90066e-315 5.50056e-315
0
9 2-In AND~
219 990 3106 0 3 22
0 22 25 111
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U24D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
6263 0 0
2
5.90066e-315 5.50185e-315
0
9 2-In AND~
219 992 3010 0 3 22
0 106 50 113
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U24C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
4900 0 0
2
5.90066e-315 5.50315e-315
0
9 2-In AND~
219 994 2902 0 3 22
0 103 26 115
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U24B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
8783 0 0
2
5.90066e-315 5.50444e-315
0
8 3-In OR~
219 1090 2891 0 4 22
0 116 115 114 108
0
0 0 608 0
4 4075
-14 -24 14 -16
4 U25A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
3221 0 0
2
5.90066e-315 5.50574e-315
0
9 2-In AND~
219 993 2948 0 3 22
0 22 26 114
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U24A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3215 0 0
2
5.90066e-315 5.50703e-315
0
9 2-In AND~
219 995 2852 0 3 22
0 106 103 116
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U23D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
7903 0 0
2
5.90066e-315 5.50833e-315
0
9 2-In AND~
219 993 2736 0 3 22
0 49 104 118
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U23C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
7121 0 0
2
5.90066e-315 5.50963e-315
0
8 3-In OR~
219 1089 2725 0 4 22
0 119 118 117 109
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
4484 0 0
2
5.90066e-315 5.51092e-315
0
9 2-In AND~
219 992 2782 0 3 22
0 22 104 117
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U23B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
5996 0 0
2
5.90066e-315 5.51222e-315
0
9 2-In AND~
219 994 2686 0 3 22
0 106 49 119
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U23A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
7804 0 0
2
5.90066e-315 5.51286e-315
0
9 2-In AND~
219 996 2525 0 3 22
0 106 102 122
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5523 0 0
2
5.90066e-315 5.51351e-315
0
9 2-In AND~
219 994 2621 0 3 22
0 22 105 120
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3330 0 0
2
5.90066e-315 5.51416e-315
0
8 3-In OR~
219 1091 2564 0 4 22
0 122 121 120 110
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
3465 0 0
2
5.90066e-315 5.51481e-315
0
9 2-In AND~
219 995 2575 0 3 22
0 102 105 121
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
8396 0 0
2
5.90066e-315 5.51545e-315
0
12 D Flip-Flop~
219 1202 2603 0 4 9
0 110 47 172 3
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U22
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3685 0 0
2
5.90066e-315 5.5161e-315
0
12 D Flip-Flop~
219 1203 2760 0 4 9
0 109 47 173 4
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U21
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7849 0 0
2
5.90066e-315 5.51675e-315
0
12 D Flip-Flop~
219 1208 3085 0 4 9
0 107 47 174 5
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U20
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6343 0 0
2
5.90066e-315 5.5174e-315
0
12 D Flip-Flop~
219 1206 2927 0 4 9
0 108 47 175 6
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U19
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7376 0 0
2
5.90066e-315 5.51804e-315
0
8 2-In OR~
219 1314 2112 0 3 22
0 124 123 102
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U18A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9156 0 0
2
5.90066e-315 5.51869e-315
0
8 4-In OR~
219 1233 2152 0 5 22
0 30 29 28 27 123
0
0 0 608 0
4 4072
-14 -24 14 -16
4 U17B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
5776 0 0
2
5.90066e-315 5.51934e-315
0
8 4-In OR~
219 1231 2073 0 5 22
0 35 34 33 32 124
0
0 0 608 0
4 4072
-14 -24 14 -16
4 U17A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
7207 0 0
2
5.90066e-315 5.51999e-315
0
9 Inverter~
13 744 2405 0 2 22
0 51 49
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U16C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
4459 0 0
2
5.90066e-315 5.52063e-315
0
9 Inverter~
13 713 2405 0 2 22
0 52 103
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U16B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
3760 0 0
2
5.90066e-315 5.52128e-315
0
9 Inverter~
13 682 2404 0 2 22
0 53 50
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U16A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
754 0 0
2
5.90066e-315 5.52193e-315
0
7 74LS154
95 1598 2840 0 22 45
0 2 2 3 4 6 5 70 71 72
73 74 75 76 77 78 79 80 81 82
83 84 85
0
0 0 4832 0
6 74F154
-21 -87 21 -79
2 U9
-7 -88 7 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
9767 0 0
2
5.90066e-315 5.52258e-315
0
5 74148
219 714 2299 0 14 29
0 2 54 55 56 57 58 59 60 61
2 53 52 51 46
0
0 0 6880 270
5 74148
-18 -60 17 -52
3 U10
56 -2 77 6
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 3 2 1 13 12 11 10
15 9 7 6 14 5 4 3 2 1
13 12 11 10 15 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
7978 0 0
2
5.90066e-315 5.52322e-315
0
14 NO PushButton~
191 195 2033 0 2 5
0 45 41
0
0 0 4704 0
0
3 S16
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3142 0 0
2
5.90066e-315 5.52387e-315
0
7 Ground~
168 238 2454 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3284 0 0
2
5.90066e-315 5.52452e-315
0
14 NO PushButton~
191 191 2243 0 2 5
0 43 41
0
0 0 4704 0
0
3 S15
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
659 0 0
2
5.90066e-315 5.52517e-315
0
14 NO PushButton~
191 194 2343 0 2 5
0 42 41
0
0 0 4704 0
0
3 S14
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3800 0 0
2
5.90066e-315 5.52581e-315
0
14 NO PushButton~
191 192 2138 0 2 5
0 44 41
0
0 0 4704 0
0
3 S13
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6792 0 0
2
5.90066e-315 5.52646e-315
0
2 +V
167 53 1977 0 1 3
0 41
0
0 0 54240 0
3 10V
-11 -23 10 -15
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3701 0 0
2
5.90066e-315 5.52711e-315
0
14 NO PushButton~
191 182 2826 0 2 5
0 39 41
0
0 0 4704 0
0
3 S12
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6316 0 0
2
5.90066e-315 5.52776e-315
0
14 NO PushButton~
191 184 3031 0 2 5
0 37 41
0
0 0 4704 0
0
3 S11
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8734 0 0
2
5.90066e-315 5.52841e-315
0
14 NO PushButton~
191 181 2931 0 2 5
0 38 41
0
0 0 4704 0
0
3 S10
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7988 0 0
2
5.90066e-315 5.52905e-315
0
7 Ground~
168 228 3142 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3217 0 0
2
5.90066e-315 5.5297e-315
0
14 NO PushButton~
191 185 2721 0 2 5
0 40 41
0
0 0 4704 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3965 0 0
2
5.90066e-315 5.53035e-315
0
14 NO PushButton~
191 1737 2047 0 2 5
0 35 36
0
0 0 4704 0
0
3 S17
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8239 0 0
2
5.90066e-315 5.531e-315
0
7 Ground~
168 1780 2468 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
828 0 0
2
5.90066e-315 5.53164e-315
0
14 NO PushButton~
191 1733 2257 0 2 5
0 33 36
0
0 0 4704 0
0
3 S18
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6187 0 0
2
5.90066e-315 5.53229e-315
0
14 NO PushButton~
191 1736 2357 0 2 5
0 32 36
0
0 0 4704 0
0
3 S19
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7107 0 0
2
5.90066e-315 5.53294e-315
0
14 NO PushButton~
191 1734 2152 0 2 5
0 34 36
0
0 0 4704 0
0
3 S20
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6433 0 0
2
5.90066e-315 5.53359e-315
0
2 +V
167 1595 1991 0 1 3
0 36
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8559 0 0
2
5.90066e-315 5.53423e-315
0
14 NO PushButton~
191 1984 2045 0 2 5
0 30 31
0
0 0 4704 0
0
3 S21
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3674 0 0
2
5.90066e-315 5.53488e-315
0
7 Ground~
168 2027 2466 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5697 0 0
2
5.90066e-315 5.53553e-315
0
14 NO PushButton~
191 1980 2255 0 2 5
0 28 31
0
0 0 4704 0
0
3 S22
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3805 0 0
2
5.90066e-315 5.53618e-315
0
14 NO PushButton~
191 1983 2355 0 2 5
0 27 31
0
0 0 4704 0
0
3 S23
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5219 0 0
2
5.90066e-315 5.53682e-315
0
14 NO PushButton~
191 1981 2150 0 2 5
0 29 31
0
0 0 4704 0
0
3 S24
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3795 0 0
2
5.90066e-315 5.53747e-315
0
2 +V
167 1842 1989 0 1 3
0 31
0
0 0 54240 0
3 15V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3637 0 0
2
5.90066e-315 5.53812e-315
0
7 Ground~
168 1209 520 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3226 0 0
2
5.90066e-315 5.53877e-315
0
5 4049~
219 1567 57 0 2 22
0 131 130
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
6966 0 0
2
5.90066e-315 5.53941e-315
0
2 +V
167 1396 71 0 1 3
0 125
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9796 0 0
2
5.90066e-315 5.54006e-315
0
14 NO PushButton~
191 1303 146 0 2 5
0 129 2
0
0 0 4704 0
0
2 S9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5952 0 0
2
5.90066e-315 5.54071e-315
0
14 NO PushButton~
191 1299 356 0 2 5
0 127 2
0
0 0 4704 0
0
2 S8
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3649 0 0
2
5.90066e-315 5.54136e-315
0
14 NO PushButton~
191 1302 456 0 2 5
0 126 2
0
0 0 4704 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3716 0 0
2
5.90066e-315 5.542e-315
0
14 NO PushButton~
191 1300 251 0 2 5
0 128 2
0
0 0 4704 0
0
2 S6
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4797 0 0
2
5.90066e-315 5.54265e-315
0
6 74LS73
102 1502 161 0 12 25
0 125 125 129 125 125 125 128 125 139
176 138 177
0
0 0 4832 0
6 74LS73
-21 -51 21 -43
3 U15
-10 -52 11 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
4681 0 0
2
5.90066e-315 5.5433e-315
0
6 74LS73
102 1503 370 0 12 25
0 125 125 127 125 125 125 126 125 137
178 136 179
0
0 0 4832 0
6 74LS73
-21 -51 21 -43
3 U14
-10 -52 11 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
9730 0 0
2
5.90066e-315 5.54395e-315
0
14 Logic Display~
6 1835 195 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9874 0 0
2
5.90066e-315 5.54459e-315
0
14 Logic Display~
6 1863 195 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
364 0 0
2
5.90066e-315 5.54524e-315
0
14 Logic Display~
6 1892 195 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3656 0 0
2
5.90066e-315 5.54589e-315
0
14 Logic Display~
6 1917 195 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3131 0 0
2
5.90066e-315 5.54654e-315
0
12 Quad D Flop~
47 1796 261 0 9 19
0 135 134 133 132 10 9 8 7 48
0
0 0 4704 0
4 QDFF
-14 -44 14 -36
3 U13
-10 -46 11 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6772 0 0
2
5.90066e-315 5.54719e-315
0
7 74LS245
64 1652 366 0 18 37
0 180 181 182 183 136 137 138 139 184
185 186 187 132 133 134 135 131 125
0
0 0 4832 0
7 74LS245
-24 -60 25 -52
3 U12
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
9557 0 0
2
5.90066e-315 5.54783e-315
0
7 74LS245
64 1665 148 0 18 37
0 188 189 190 191 105 104 26 25 192
193 194 195 132 133 134 135 130 125
0
0 0 4832 0
7 74LS245
-24 -60 25 -52
3 U11
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
5789 0 0
2
5.90066e-315 5.54848e-315
0
5 4049~
219 272 1033 0 2 22
0 141 140
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
7328 0 0
2
44974.9 21
0
14 NO PushButton~
191 213 1131 0 2 5
0 142 143
0
0 0 4704 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4799 0 0
2
44974.9 22
0
14 Logic Display~
6 813 1277 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9196 0 0
2
44974.9 23
0
14 Logic Display~
6 812 1190 0 1 2
10 131
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3857 0 0
2
44974.9 24
0
14 Logic Display~
6 815 1093 0 1 2
10 144
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7125 0 0
2
44974.9 25
0
4 4017
219 552 1165 0 14 29
0 140 142 145 22 131 144 145 196 197
198 199 200 201 202
0
0 0 6880 0
4 4017
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
3641 0 0
2
44974.9 26
0
5 4049~
219 278 475 0 2 22
0 152 147
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
9821 0 0
2
44974.9 27
0
14 NO PushButton~
191 229 871 0 2 5
0 149 143
0
0 0 4704 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3187 0 0
2
44974.9 28
0
5 4049~
219 229 527 0 2 22
0 149 150
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
762 0 0
2
44974.9 29
0
9 2-In AND~
219 240 567 0 3 22
0 150 13 151
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
39 0 0
2
44974.9 30
0
14 Logic Display~
6 815 1032 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9450 0 0
2
44974.9 31
0
14 Logic Display~
6 817 957 0 1 2
10 141
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3236 0 0
2
44974.9 32
0
14 Logic Display~
6 816 904 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3321 0 0
2
5.90066e-315 5.54913e-315
0
9 2-In AND~
219 771 924 0 3 22
0 146 152 48
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8879 0 0
2
5.90066e-315 5.54978e-315
0
14 NO PushButton~
191 229 834 0 2 5
0 153 143
0
0 0 4704 0
0
2 S2
-7 -22 7 -14
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5433 0 0
2
5.90066e-315 5.55042e-315
0
5 4049~
219 202 386 0 2 22
0 153 155
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
3679 0 0
2
5.90066e-315 5.55107e-315
0
9 2-In AND~
219 224 427 0 3 22
0 155 146 154
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9342 0 0
2
5.90066e-315 5.55172e-315
0
5 4049~
219 190 297 0 2 22
0 158 157
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3623 0 0
2
5.90066e-315 5.55237e-315
0
7 Ground~
168 357 1484 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3722 0 0
2
5.90066e-315 5.55301e-315
0
2 +V
167 163 761 0 1 3
0 143
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8993 0 0
2
5.90066e-315 5.55366e-315
0
14 NO PushButton~
191 227 794 0 2 5
0 158 143
0
0 0 4704 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3723 0 0
2
5.90066e-315 5.55398e-315
0
8 3-In OR~
219 299 352 0 4 22
0 156 151 154 159
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
6244 0 0
2
5.90066e-315 5.55431e-315
0
9 2-In AND~
219 220 350 0 3 22
0 157 141 156
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6421 0 0
2
5.90066e-315 5.55463e-315
0
7 Ground~
168 864 600 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7743 0 0
2
5.90066e-315 5.55496e-315
0
4 LED~
171 949 545 0 2 2
10 160 2
0
0 0 864 0
4 LED1
17 0 45 8
3 D13
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9840 0 0
2
5.90066e-315 5.55528e-315
0
4 LED~
171 908 540 0 2 2
10 161 2
0
0 0 864 0
4 LED1
17 0 45 8
3 D12
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6910 0 0
2
5.90066e-315 5.5556e-315
0
4 LED~
171 856 539 0 2 2
10 162 2
0
0 0 864 0
4 LED1
17 0 45 8
3 D11
20 -10 41 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
449 0 0
2
5.90066e-315 5.55593e-315
0
4 LED~
171 802 541 0 2 2
10 148 2
0
0 0 864 0
4 LED1
17 0 45 8
3 D10
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8761 0 0
2
5.90066e-315 5.55625e-315
0
4 LED~
171 744 535 0 2 2
10 13 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D9
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6748 0 0
2
5.90066e-315 5.55657e-315
0
4 LED~
171 685 535 0 2 2
10 146 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7393 0 0
2
5.90066e-315 5.5569e-315
0
4 LED~
171 625 534 0 2 2
10 141 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7699 0 0
2
5.90066e-315 5.55722e-315
0
4 LED~
171 568 532 0 2 2
10 163 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6638 0 0
2
5.90066e-315 5.55755e-315
0
4 LED~
171 509 531 0 2 2
10 164 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4595 0 0
2
5.90066e-315 5.55787e-315
0
4 4017
219 434 448 0 14 29
0 159 147 148 164 163 141 146 13 148
162 161 160 165 203
0
0 0 6880 0
4 4017
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
9395 0 0
2
5.90066e-315 5.55819e-315
0
7 Ground~
168 940 271 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3303 0 0
2
5.90066e-315 5.55852e-315
0
7 Pulser~
4 40 35 0 10 12
0 204 205 152 206 0 0 5 5 4
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4498 0 0
2
5.90066e-315 5.55884e-315
0
9 2-In AND~
219 192 163 0 3 22
0 152 163 167
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9728 0 0
2
44974.9 33
0
4 LED~
171 895 231 0 2 2
10 25 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3789 0 0
2
44974.9 34
0
4 LED~
171 834 229 0 2 2
10 26 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3978 0 0
2
44974.9 35
0
4 LED~
171 776 227 0 2 2
10 104 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3494 0 0
2
44974.9 36
0
4 LED~
171 716 223 0 2 2
10 105 2
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3507 0 0
2
44974.9 37
0
7 74LS175
131 652 147 0 14 29
0 171 167 170 169 168 166 105 207 104
208 26 209 25 210
0
0 0 4832 0
7 74LS175
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 9 13 12 5 4 15 14 10
11 7 6 2 3 1 9 13 12 5
4 15 14 10 11 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
5151 0 0
2
44974.9 38
0
2 +V
167 503 30 0 1 3
0 171
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3701 0 0
2
44974.9 39
0
7 Ground~
168 268 194 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8585 0 0
2
44974.9 40
0
7 74LS161
96 377 86 0 14 29
0 171 171 152 2 2 2 2 171 171
211 166 168 169 170
0
0 0 6880 0
8 74LS161A
-28 -60 28 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
8809 0 0
2
44974.9 41
0
9 Resistor~
219 238 2402 0 3 5
0 2 42 -1
0
0 0 864 90
2 1k
8 0 22 8
3 R16
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5993 0 0
2
5.90066e-315 5.55917e-315
0
9 Resistor~
219 111 2272 0 4 5
0 43 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R15
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8654 0 0
2
5.90066e-315 5.55949e-315
0
9 Resistor~
219 110 2166 0 4 5
0 44 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R14
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7223 0 0
2
5.90066e-315 5.55981e-315
0
9 Resistor~
219 109 2061 0 4 5
0 45 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3641 0 0
2
5.90066e-315 5.56014e-315
0
9 Resistor~
219 99 2749 0 4 5
0 40 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3104 0 0
2
5.90066e-315 5.56046e-315
0
9 Resistor~
219 100 2854 0 4 5
0 39 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3296 0 0
2
5.90066e-315 5.56078e-315
0
9 Resistor~
219 101 2960 0 4 5
0 38 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8534 0 0
2
5.90066e-315 5.56111e-315
0
9 Resistor~
219 228 3090 0 3 5
0 2 37 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
949 0 0
2
5.90066e-315 5.56143e-315
0
9 Resistor~
219 1780 2416 0 3 5
0 2 32 -1
0
0 0 864 90
2 1k
11 0 25 8
3 R17
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3371 0 0
2
5.90066e-315 5.56176e-315
0
9 Resistor~
219 1653 2286 0 4 5
0 33 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R18
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7311 0 0
2
5.90066e-315 5.56208e-315
0
9 Resistor~
219 1652 2180 0 4 5
0 34 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R19
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
5.90066e-315 5.5624e-315
0
9 Resistor~
219 1651 2075 0 4 5
0 35 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R20
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3526 0 0
2
5.90066e-315 5.56273e-315
0
9 Resistor~
219 2027 2414 0 3 5
0 2 27 -1
0
0 0 864 90
2 1k
11 0 25 8
3 R21
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4129 0 0
2
5.90066e-315 5.56305e-315
0
9 Resistor~
219 1900 2284 0 4 5
0 28 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R22
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6278 0 0
2
5.90066e-315 5.56337e-315
0
9 Resistor~
219 1899 2178 0 4 5
0 29 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R23
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3482 0 0
2
5.90066e-315 5.5637e-315
0
9 Resistor~
219 1898 2073 0 4 5
0 30 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R24
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8323 0 0
2
5.90066e-315 5.56402e-315
0
9 Resistor~
219 1355 440 0 4 5
0 126 125 0 1
0
0 0 864 0
2 1k
-7 -15 7 -7
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3984 0 0
2
5.90066e-315 5.56435e-315
0
9 Resistor~
219 1348 336 0 4 5
0 127 125 0 1
0
0 0 864 0
2 1k
-7 -15 7 -7
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7622 0 0
2
5.90066e-315 5.56467e-315
0
9 Resistor~
219 1335 220 0 4 5
0 128 125 0 1
0
0 0 864 0
2 1k
-7 -15 7 -7
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
816 0 0
2
5.90066e-315 5.56499e-315
0
9 Resistor~
219 1347 117 0 4 5
0 129 125 0 1
0
0 0 864 0
2 1k
-7 -15 7 -7
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4656 0 0
2
5.90066e-315 5.56532e-315
0
9 Resistor~
219 275 1140 0 4 5
0 142 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R2
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6356 0 0
2
44974.9 42
0
9 Resistor~
219 282 879 0 4 5
0 149 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R4
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7479 0 0
2
44974.9 43
0
9 Resistor~
219 280 841 0 4 5
0 153 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R3
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5690 0 0
2
5.90066e-315 5.56564e-315
0
9 Resistor~
219 275 803 0 4 5
0 158 2 0 -1
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R1
-9 -24 5 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5617 0 0
2
44974.9 44
0
420
0 0 3 0 0 8320 0 0 0 30 211 5
2233 1396
2501 1396
2501 2997
1521 2997
1521 2858
0 0 4 0 0 12416 0 0 0 210 31 5
1512 2867
1512 3008
2512 3008
2512 1388
2188 1388
0 0 5 0 0 12416 0 0 0 208 33 5
1496 2885
1496 3024
2533 3024
2533 1363
2099 1363
0 0 6 0 0 16512 0 0 0 32 209 7
2150 1376
2553 1376
2553 1713
2521 1713
2521 3012
1503 3012
1503 2876
0 0 7 0 0 8320 0 0 0 34 288 5
2023 1397
1839 1397
1839 324
1886 324
1886 267
0 0 8 0 0 4224 0 0 0 289 35 3
1858 255
1858 1390
1982 1390
0 0 9 0 0 8320 0 0 0 36 290 5
1943 1377
1930 1377
1930 300
1841 300
1841 243
5 0 10 0 0 4224 0 140 0 0 37 3
1820 231
1820 1368
1901 1368
3 1 11 0 0 8320 0 18 21 0 0 5
2698 1572
2712 1572
2712 1619
2759 1619
2759 1586
3 1 12 0 0 8320 0 17 20 0 0 5
2697 1403
2712 1403
2712 1463
2764 1463
2764 1416
1 1 13 0 0 16384 0 17 18 0 0 6
2652 1394
2616 1394
2616 1349
2638 1349
2638 1563
2653 1563
1 0 13 0 0 0 0 19 0 0 11 5
2669 1286
2711 1286
2711 1348
2638 1348
2638 1349
2 2 14 0 0 4224 0 16 17 0 0 3
2616 1451
2616 1412
2652 1412
3 2 15 0 0 12416 0 15 18 0 0 4
2515 1509
2568 1509
2568 1581
2653 1581
3 1 15 0 0 0 0 15 16 0 0 4
2515 1509
2568 1509
2568 1451
2580 1451
3 2 16 0 0 4224 0 14 15 0 0 3
2430 1567
2430 1518
2469 1518
3 1 17 0 0 4224 0 13 15 0 0 3
2435 1451
2435 1500
2469 1500
3 2 18 0 0 8320 0 12 14 0 0 3
2342 1609
2342 1576
2384 1576
3 1 19 0 0 8320 0 11 14 0 0 3
2339 1544
2339 1558
2384 1558
3 2 20 0 0 8320 0 10 13 0 0 3
2339 1480
2339 1460
2389 1460
3 1 21 0 0 8320 0 9 13 0 0 3
2340 1418
2340 1442
2389 1442
2 0 3 0 0 0 0 12 0 0 30 2
2293 1618
2233 1618
1 0 7 0 0 0 0 12 0 0 34 2
2293 1600
2023 1600
2 0 4 0 0 0 0 11 0 0 31 2
2290 1553
2188 1553
1 0 8 0 0 0 0 11 0 0 35 2
2290 1535
1982 1535
2 0 6 0 0 0 0 10 0 0 32 2
2290 1489
2150 1489
1 0 9 0 0 0 0 10 0 0 36 2
2290 1471
1943 1471
2 0 5 0 0 0 0 9 0 0 33 2
2291 1427
2099 1427
1 0 10 0 0 0 0 9 0 0 37 2
2291 1409
1901 1409
0 0 3 0 0 0 0 0 0 38 0 3
2254 1346
2233 1346
2233 1752
0 0 4 0 0 0 0 0 0 40 0 3
2210 1344
2188 1344
2188 1749
0 0 6 0 0 0 0 0 0 42 0 3
2168 1345
2150 1345
2150 1754
0 0 5 0 0 0 0 0 0 44 0 3
2124 1343
2099 1343
2099 1751
0 0 7 0 0 0 0 0 0 46 0 3
2045 1344
2023 1344
2023 1755
0 0 8 0 0 0 0 0 0 48 0 3
2005 1345
1982 1345
1982 1753
0 0 9 0 0 0 0 0 0 50 0 3
1961 1343
1943 1343
1943 1755
0 0 10 0 0 0 0 0 0 52 0 3
1920 1344
1901 1344
1901 1754
1 0 3 0 0 0 0 1 0 0 39 2
2254 1324
2254 1346
0 1 3 0 0 0 0 0 1 0 0 2
2254 1350
2254 1324
1 0 4 0 0 0 0 2 0 0 41 2
2210 1323
2210 1345
0 1 4 0 0 0 0 0 2 0 0 2
2210 1349
2210 1323
1 0 6 0 0 0 0 3 0 0 43 2
2168 1323
2168 1345
0 1 6 0 0 0 0 0 3 0 0 2
2168 1349
2168 1323
1 0 5 0 0 0 0 4 0 0 45 2
2124 1322
2124 1344
0 1 5 0 0 0 0 0 4 0 0 2
2124 1348
2124 1322
1 0 7 0 0 0 0 5 0 0 47 2
2045 1323
2045 1345
0 1 7 0 0 0 0 0 5 0 0 2
2045 1349
2045 1323
1 0 8 0 0 0 0 6 0 0 49 2
2005 1323
2005 1345
0 1 8 0 0 0 0 0 6 0 0 2
2005 1349
2005 1323
1 0 9 0 0 0 0 7 0 0 51 2
1961 1322
1961 1344
0 1 9 0 0 0 0 0 7 0 0 2
1961 1348
1961 1322
1 0 10 0 0 0 0 8 0 0 53 2
1920 1322
1920 1344
0 1 10 0 0 0 0 0 8 0 0 2
1920 1348
1920 1322
2 0 22 0 0 4096 0 22 0 0 315 2
1081 2439
549 2439
1 2 23 0 0 4224 0 22 23 0 0 4
1081 2421
908 2421
908 2372
866 2372
3 1 24 0 0 8320 0 22 24 0 0 6
1127 2430
1150 2430
1150 2774
1196 2774
1196 2795
1200 2795
2 0 2 0 0 4096 0 197 0 0 97 2
1635 2286
1620 2286
1 0 22 0 0 0 0 75 0 0 315 3
522 3156
522 3170
538 3170
0 0 25 0 0 4096 0 0 0 402 0 2
994 174
1137 174
0 0 26 0 0 4096 0 0 0 403 0 2
983 156
1138 156
0 0 2 0 0 12288 0 0 0 175 97 5
1507 2748
1507 2714
1752 2714
1752 2454
1780 2454
0 4 27 0 0 8192 0 0 97 71 0 7
2014 2363
2014 2168
1275 2168
1275 2177
1183 2177
1183 2166
1216 2166
0 3 28 0 0 8192 0 0 97 73 0 5
1960 2284
1960 2273
1188 2273
1188 2157
1216 2157
0 2 29 0 0 8192 0 0 97 69 0 7
1967 2178
1967 2168
1270 2168
1270 2172
1193 2172
1193 2148
1216 2148
0 1 30 0 0 8192 0 0 97 78 0 5
1966 2073
1966 2132
1193 2132
1193 2139
1216 2139
0 1 27 0 0 12416 0 0 34 71 0 5
2027 2363
2021 2363
2021 2014
1107 2014
1107 2029
0 1 29 0 0 8320 0 0 36 69 0 4
2006 2158
2006 2010
958 2010
958 2025
0 1 30 0 0 12416 0 0 37 78 0 5
2009 2054
2005 2054
2005 2005
901 2005
901 2025
1 1 29 0 0 0 0 202 125 0 0 4
1917 2178
2006 2178
2006 2158
1998 2158
0 2 31 0 0 4096 0 0 125 82 0 2
1842 2158
1964 2158
2 1 27 0 0 0 0 200 124 0 0 3
2027 2396
2027 2363
2000 2363
0 2 31 0 0 4096 0 0 124 82 0 3
1842 2361
1966 2361
1966 2363
1 1 28 0 0 0 0 123 201 0 0 4
1997 2263
2001 2263
2001 2284
1918 2284
0 2 31 0 0 0 0 0 123 82 0 2
1842 2263
1963 2263
1 1 28 0 0 8320 0 35 123 0 0 5
1042 2026
1042 2006
2015 2006
2015 2263
1997 2263
1 2 2 0 0 12288 0 122 203 0 0 5
2027 2460
2027 2436
1867 2436
1867 2073
1880 2073
1 1 2 0 0 0 0 122 200 0 0 2
2027 2460
2027 2432
1 1 30 0 0 0 0 203 121 0 0 4
1916 2073
2009 2073
2009 2053
2001 2053
0 2 31 0 0 4096 0 0 121 82 0 2
1842 2053
1967 2053
0 2 2 0 0 0 0 0 202 76 0 4
1867 2179
1871 2179
1871 2178
1881 2178
0 2 2 0 0 0 0 0 201 76 0 4
1867 2286
1871 2286
1871 2284
1882 2284
1 0 31 0 0 4224 0 126 0 0 0 2
1842 1998
1842 2648
4 0 32 0 0 12288 0 98 0 0 92 4
1214 2087
1200 2087
1200 2390
1780 2390
3 0 33 0 0 12288 0 98 0 0 94 5
1214 2078
1205 2078
1205 2295
1713 2295
1713 2286
2 0 34 0 0 12288 0 98 0 0 90 5
1214 2069
1210 2069
1210 2189
1716 2189
1716 2180
1 0 35 0 0 12288 0 98 0 0 99 5
1214 2060
1210 2060
1210 2033
1715 2033
1715 2075
0 1 32 0 0 12416 0 0 38 92 0 5
1780 2367
1774 2367
1774 2007
818 2007
818 2027
0 1 34 0 0 8320 0 0 40 90 0 4
1759 2160
1759 2004
674 2004
674 2029
0 1 35 0 0 12416 0 0 41 99 0 5
1762 2057
1758 2057
1758 2004
612 2004
612 2031
1 1 34 0 0 0 0 198 119 0 0 4
1670 2180
1759 2180
1759 2160
1751 2160
0 2 36 0 0 4096 0 0 119 103 0 2
1595 2160
1717 2160
2 1 32 0 0 0 0 196 118 0 0 3
1780 2398
1780 2365
1753 2365
0 2 36 0 0 4096 0 0 118 103 0 2
1595 2365
1719 2365
1 1 33 0 0 0 0 117 197 0 0 4
1750 2265
1754 2265
1754 2286
1671 2286
0 2 36 0 0 0 0 0 117 103 0 2
1595 2265
1716 2265
1 1 33 0 0 8320 0 39 117 0 0 5
755 2029
755 2004
1768 2004
1768 2265
1750 2265
1 2 2 0 0 0 0 116 199 0 0 5
1780 2462
1780 2438
1620 2438
1620 2075
1633 2075
1 1 2 0 0 0 0 116 196 0 0 2
1780 2462
1780 2434
1 1 35 0 0 0 0 199 115 0 0 4
1669 2075
1762 2075
1762 2055
1754 2055
0 2 36 0 0 4096 0 0 115 103 0 2
1595 2055
1720 2055
0 2 2 0 0 0 0 0 198 97 0 2
1620 2180
1634 2180
0 2 2 0 0 0 0 0 197 0 0 2
1624 2286
1635 2286
1 0 36 0 0 4224 0 120 0 0 0 2
1595 2000
1595 2650
2 0 37 0 0 12416 0 34 0 0 120 5
1089 2029
1089 1958
362 1958
362 3039
228 3039
2 0 38 0 0 12416 0 35 0 0 114 6
1024 2026
1024 1998
217 1998
217 2934
212 2934
212 2939
0 2 39 0 0 8320 0 0 36 117 0 5
213 2834
931 2834
931 2010
940 2010
940 2025
0 2 40 0 0 8320 0 0 37 115 0 5
214 2731
875 2731
875 2010
883 2010
883 2025
1 1 38 0 0 0 0 112 194 0 0 4
198 2939
202 2939
202 2960
119 2960
2 0 41 0 0 4096 0 111 0 0 113 2
167 3039
45 3039
2 0 41 0 0 0 0 112 0 0 113 2
164 2939
45 2939
2 0 41 0 0 4096 0 114 0 0 113 2
168 2729
45 2729
2 0 41 0 0 0 0 110 0 0 113 2
165 2834
45 2834
0 0 41 0 0 8192 0 0 0 131 0 3
47 2674
45 2674
45 3324
1 0 38 0 0 0 0 112 0 0 0 2
198 2939
216 2939
1 1 40 0 0 0 0 192 114 0 0 4
117 2749
214 2749
214 2729
202 2729
2 1 2 0 0 8192 0 192 113 0 0 5
81 2749
72 2749
72 3127
228 3127
228 3136
1 1 39 0 0 0 0 193 110 0 0 4
118 2854
213 2854
213 2834
199 2834
2 0 2 0 0 0 0 193 0 0 116 2
82 2854
72 2854
2 0 2 0 0 0 0 194 0 0 116 2
83 2960
72 2960
2 1 37 0 0 0 0 195 111 0 0 3
228 3072
228 3039
201 3039
1 1 2 0 0 0 0 113 195 0 0 2
228 3136
228 3108
0 2 42 0 0 4224 0 0 38 138 0 5
238 2352
793 2352
793 2012
800 2012
800 2027
0 2 43 0 0 8320 0 0 39 132 0 4
221 2251
221 2004
737 2004
737 2029
0 2 44 0 0 4224 0 0 40 135 0 5
223 2146
585 2146
585 2009
656 2009
656 2029
0 2 45 0 0 4224 0 0 41 133 0 5
224 2041
591 2041
591 2016
594 2016
594 2031
1 1 43 0 0 0 0 106 189 0 0 4
208 2251
212 2251
212 2272
129 2272
2 0 41 0 0 0 0 107 0 0 131 2
177 2351
47 2351
2 0 41 0 0 0 0 106 0 0 131 2
174 2251
47 2251
2 0 41 0 0 0 0 104 0 0 131 2
178 2041
47 2041
2 0 41 0 0 0 0 108 0 0 131 2
175 2146
47 2146
1 0 41 0 0 8320 0 109 0 0 113 4
53 1986
47 1986
47 2679
45 2679
1 0 43 0 0 0 0 106 0 0 0 2
208 2251
226 2251
1 1 45 0 0 0 0 191 104 0 0 4
127 2061
224 2061
224 2041
212 2041
2 1 2 0 0 0 0 191 105 0 0 5
91 2061
82 2061
82 2439
238 2439
238 2448
1 1 44 0 0 0 0 190 108 0 0 4
128 2166
223 2166
223 2146
209 2146
2 0 2 0 0 0 0 190 0 0 134 2
92 2166
82 2166
2 0 2 0 0 0 0 189 0 0 134 2
93 2272
82 2272
2 1 42 0 0 0 0 188 107 0 0 3
238 2384
238 2351
211 2351
1 1 2 0 0 0 0 105 188 0 0 2
238 2448
238 2420
14 1 46 0 0 8320 0 103 23 0 0 3
752 2339
752 2372
830 2372
3 2 47 0 0 8320 0 24 94 0 0 6
1245 2804
1259 2804
1259 3082
1176 3082
1176 3067
1184 3067
3 2 47 0 0 0 0 24 95 0 0 6
1245 2804
1248 2804
1248 2924
1174 2924
1174 2909
1182 2909
0 2 47 0 0 0 0 0 92 144 0 5
1249 2804
1249 2600
1170 2600
1170 2585
1178 2585
3 2 47 0 0 0 0 24 93 0 0 6
1245 2804
1249 2804
1249 2757
1166 2757
1166 2742
1179 2742
0 2 48 0 0 12416 0 0 24 287 0 9
1469 924
1469 1426
409 1426
409 2817
1071 2817
1071 2790
1157 2790
1157 2813
1200 2813
1 0 49 0 0 4096 0 84 0 0 147 3
969 2727
920 2727
920 2695
2 2 49 0 0 4224 0 99 87 0 0 3
747 2423
747 2695
970 2695
1 0 50 0 0 4096 0 76 0 0 149 3
967 3051
930 3051
930 3019
2 2 50 0 0 4224 0 101 79 0 0 3
685 2422
685 3019
968 3019
1 0 22 0 0 0 0 78 0 0 315 2
966 3097
549 3097
1 0 22 0 0 0 0 82 0 0 315 2
969 2939
549 2939
1 0 22 0 0 0 0 86 0 0 315 2
968 2773
549 2773
1 0 22 0 0 0 0 89 0 0 315 2
970 2612
549 2612
1 1 2 0 0 0 0 103 25 0 0 4
752 2263
752 2259
824 2259
824 2291
13 1 51 0 0 4224 0 103 99 0 0 4
725 2339
725 2379
747 2379
747 2387
12 1 52 0 0 4224 0 103 100 0 0 2
716 2339
716 2387
11 1 53 0 0 4224 0 103 101 0 0 4
707 2339
707 2378
685 2378
685 2386
2 2 54 0 0 8320 0 26 103 0 0 4
1098 2150
1098 2231
734 2231
734 2263
2 3 55 0 0 8320 0 27 103 0 0 4
1033 2151
1033 2236
725 2236
725 2263
2 4 56 0 0 8320 0 28 103 0 0 4
953 2151
953 2241
716 2241
716 2263
2 5 57 0 0 8320 0 29 103 0 0 4
890 2150
890 2246
707 2246
707 2263
2 6 58 0 0 8320 0 30 103 0 0 4
808 2150
808 2250
698 2250
698 2263
2 7 59 0 0 4224 0 31 103 0 0 4
747 2151
747 2255
689 2255
689 2263
2 8 60 0 0 4224 0 32 103 0 0 4
663 2149
663 2250
680 2250
680 2263
2 9 61 0 0 4224 0 33 103 0 0 4
606 2150
606 2255
671 2255
671 2263
3 1 62 0 0 4224 0 34 26 0 0 2
1098 2075
1098 2114
3 1 63 0 0 4224 0 35 27 0 0 2
1033 2072
1033 2115
3 1 64 0 0 4224 0 36 28 0 0 4
949 2071
949 2107
953 2107
953 2115
3 1 65 0 0 4224 0 37 29 0 0 4
892 2071
892 2106
890 2106
890 2114
3 1 66 0 0 4224 0 38 30 0 0 4
809 2073
809 2106
808 2106
808 2114
3 1 67 0 0 4224 0 39 31 0 0 4
746 2075
746 2107
747 2107
747 2115
3 1 68 0 0 4224 0 40 32 0 0 4
665 2075
665 2105
663 2105
663 2113
3 1 69 0 0 4224 0 41 33 0 0 4
603 2077
603 2106
606 2106
606 2114
10 1 2 0 0 0 0 103 42 0 0 6
671 2339
671 2347
640 2347
640 2312
623 2312
623 2326
2 1 2 0 0 0 0 102 102 0 0 8
1560 2831
1518 2831
1518 2785
1488 2785
1488 2748
1531 2748
1531 2822
1560 2822
7 1 70 0 0 4224 0 102 46 0 0 3
1636 2777
2479 2777
2479 2655
8 1 71 0 0 4224 0 102 45 0 0 3
1636 2786
2446 2786
2446 2656
9 1 72 0 0 4224 0 102 44 0 0 3
1636 2795
2414 2795
2414 2655
10 1 73 0 0 4224 0 102 43 0 0 3
1636 2804
2379 2804
2379 2659
11 1 74 0 0 4224 0 102 50 0 0 3
1636 2813
2310 2813
2310 2655
12 1 75 0 0 4224 0 102 49 0 0 3
1636 2822
2277 2822
2277 2656
13 1 76 0 0 4224 0 102 48 0 0 3
1636 2831
2245 2831
2245 2655
14 1 77 0 0 4224 0 102 47 0 0 3
1636 2840
2210 2840
2210 2659
15 1 78 0 0 4224 0 102 54 0 0 3
1636 2849
2141 2849
2141 2656
16 1 79 0 0 4224 0 102 53 0 0 3
1636 2858
2108 2858
2108 2657
17 1 80 0 0 4224 0 102 52 0 0 3
1636 2867
2076 2867
2076 2656
18 1 81 0 0 4224 0 102 51 0 0 3
1636 2876
2041 2876
2041 2660
19 1 82 0 0 4224 0 102 55 0 0 3
1636 2885
1977 2885
1977 2660
20 1 83 0 0 4224 0 102 56 0 0 3
1636 2894
1944 2894
1944 2661
21 1 84 0 0 4224 0 102 57 0 0 3
1636 2903
1912 2903
1912 2660
22 1 85 0 0 8320 0 102 74 0 0 3
1636 2912
1877 2912
1877 2664
1 2 86 0 0 8320 0 69 46 0 0 3
2478 2610
2479 2610
2479 2619
1 2 87 0 0 8320 0 70 45 0 0 3
2445 2609
2446 2609
2446 2620
1 2 88 0 0 8320 0 71 44 0 0 3
2413 2609
2414 2609
2414 2619
1 2 89 0 0 8320 0 72 43 0 0 3
2378 2610
2379 2610
2379 2623
1 2 90 0 0 8320 0 65 50 0 0 3
2309 2610
2310 2610
2310 2619
1 2 91 0 0 8320 0 66 49 0 0 3
2276 2609
2277 2609
2277 2620
1 2 92 0 0 8320 0 67 48 0 0 3
2244 2609
2245 2609
2245 2619
1 2 93 0 0 8320 0 68 47 0 0 3
2209 2610
2210 2610
2210 2623
1 2 94 0 0 4224 0 62 54 0 0 2
2141 2611
2141 2620
1 2 95 0 0 4224 0 73 53 0 0 2
2108 2610
2108 2621
1 2 96 0 0 4224 0 63 52 0 0 2
2076 2610
2076 2620
1 2 97 0 0 4224 0 64 51 0 0 2
2041 2611
2041 2624
1 2 98 0 0 4224 0 61 55 0 0 2
1977 2613
1977 2624
1 2 99 0 0 4224 0 60 56 0 0 2
1944 2612
1944 2625
1 2 100 0 0 4224 0 59 57 0 0 2
1912 2612
1912 2624
1 2 101 0 0 4224 0 58 74 0 0 2
1877 2613
1877 2628
4 6 5 0 0 0 0 94 102 0 0 4
1232 3049
1409 3049
1409 2885
1566 2885
4 5 6 0 0 0 0 95 102 0 0 4
1230 2891
1386 2891
1386 2876
1566 2876
4 4 4 0 0 0 0 93 102 0 0 4
1227 2724
1385 2724
1385 2867
1566 2867
4 3 3 0 0 0 0 92 102 0 0 4
1226 2567
1409 2567
1409 2858
1566 2858
1 0 102 0 0 8192 0 91 0 0 223 3
971 2566
949 2566
949 2534
1 0 103 0 0 4096 0 80 0 0 214 3
970 2893
930 2893
930 2861
2 2 103 0 0 4224 0 100 83 0 0 3
716 2423
716 2861
971 2861
2 0 25 0 0 4096 0 78 0 0 245 2
966 3115
808 3115
2 0 25 0 0 4096 0 76 0 0 245 2
967 3069
808 3069
2 0 26 0 0 4096 0 82 0 0 246 2
969 2957
737 2957
2 0 26 0 0 4096 0 80 0 0 246 2
970 2911
737 2911
2 0 104 0 0 4096 0 86 0 0 247 2
968 2791
674 2791
2 0 104 0 0 4096 0 84 0 0 247 2
969 2745
674 2745
2 0 105 0 0 4096 0 89 0 0 248 2
970 2630
612 2630
2 0 105 0 0 4096 0 91 0 0 248 2
971 2584
612 2584
3 2 102 0 0 12416 0 96 88 0 0 6
1347 2112
1424 2112
1424 2358
934 2358
934 2534
972 2534
1 0 106 0 0 4096 0 79 0 0 228 2
968 3001
522 3001
1 0 106 0 0 4096 0 83 0 0 228 2
971 2843
522 2843
1 0 106 0 0 0 0 87 0 0 228 2
970 2677
522 2677
1 0 106 0 0 4096 0 88 0 0 228 2
972 2516
522 2516
2 0 106 0 0 4224 0 75 0 0 0 2
522 3120
522 2422
4 1 107 0 0 4224 0 77 94 0 0 2
1120 3049
1184 3049
4 1 108 0 0 4224 0 81 95 0 0 2
1123 2891
1182 2891
4 1 109 0 0 8320 0 85 93 0 0 3
1122 2725
1122 2724
1179 2724
4 1 110 0 0 8320 0 90 92 0 0 3
1124 2564
1124 2567
1178 2567
3 3 111 0 0 4224 0 78 77 0 0 4
1011 3106
1068 3106
1068 3058
1074 3058
3 2 112 0 0 4224 0 76 77 0 0 4
1012 3060
1056 3060
1056 3049
1075 3049
3 1 113 0 0 4224 0 79 77 0 0 4
1013 3010
1051 3010
1051 3040
1074 3040
3 3 114 0 0 4224 0 82 81 0 0 4
1014 2948
1071 2948
1071 2900
1077 2900
3 2 115 0 0 4224 0 80 81 0 0 4
1015 2902
1059 2902
1059 2891
1078 2891
3 1 116 0 0 4224 0 83 81 0 0 4
1016 2852
1054 2852
1054 2882
1077 2882
3 3 117 0 0 4224 0 86 85 0 0 4
1013 2782
1070 2782
1070 2734
1076 2734
3 2 118 0 0 4224 0 84 85 0 0 4
1014 2736
1058 2736
1058 2725
1077 2725
3 1 119 0 0 4224 0 87 85 0 0 4
1015 2686
1053 2686
1053 2716
1076 2716
3 3 120 0 0 4224 0 89 90 0 0 4
1015 2621
1072 2621
1072 2573
1078 2573
3 2 121 0 0 4224 0 91 90 0 0 4
1016 2575
1060 2575
1060 2564
1079 2564
3 1 122 0 0 4224 0 88 90 0 0 4
1017 2525
1055 2525
1055 2555
1078 2555
0 0 25 0 0 12416 0 0 0 59 0 6
1012 174
1012 1538
33 1538
33 3297
808 3297
808 2503
0 0 26 0 0 12416 0 0 0 60 0 6
1048 156
1048 1504
7 1504
7 3284
737 3284
737 2503
0 0 104 0 0 12416 0 0 0 404 0 6
1039 138
1039 1514
16 1514
16 3259
674 3259
674 2502
0 0 105 0 0 12416 0 0 0 405 0 6
1023 120
1023 1527
23 1527
23 3269
612 3269
612 2420
5 2 123 0 0 8320 0 97 96 0 0 4
1266 2152
1277 2152
1277 2121
1301 2121
5 1 124 0 0 8320 0 98 96 0 0 4
1264 2073
1277 2073
1277 2103
1301 2103
0 18 125 0 0 4096 0 0 142 305 0 4
1396 244
1731 244
1731 112
1697 112
2 0 125 0 0 0 0 204 0 0 305 2
1373 440
1396 440
2 0 125 0 0 0 0 205 0 0 305 2
1366 336
1396 336
2 0 125 0 0 0 0 206 0 0 305 2
1353 220
1396 220
2 0 125 0 0 0 0 207 0 0 305 2
1365 117
1396 117
1 0 126 0 0 4096 0 204 0 0 294 2
1337 440
1337 463
1 0 127 0 0 4096 0 205 0 0 292 2
1330 336
1330 364
1 1 128 0 0 4096 0 206 133 0 0 2
1317 220
1317 259
1 0 129 0 0 4096 0 207 0 0 264 2
1329 117
1329 152
2 0 2 0 0 0 0 132 0 0 266 2
1285 464
1209 464
2 0 2 0 0 0 0 131 0 0 266 2
1282 364
1209 364
1 7 128 0 0 12416 0 133 134 0 0 4
1317 259
1363 259
1363 188
1464 188
2 0 2 0 0 0 0 133 0 0 266 2
1283 259
1209 259
1 3 129 0 0 8320 0 130 134 0 0 3
1320 154
1320 152
1464 152
2 0 2 0 0 0 0 130 0 0 266 2
1286 154
1209 154
0 1 2 0 0 4096 0 0 127 0 0 2
1209 71
1209 514
8 0 125 0 0 0 0 134 0 0 305 2
1464 197
1396 197
5 0 105 0 0 0 0 142 0 0 405 5
1633 157
1614 157
1614 41
893 41
893 120
6 0 104 0 0 0 0 142 0 0 404 5
1633 166
1608 166
1608 30
912 30
912 138
7 0 26 0 0 0 0 142 0 0 403 5
1633 175
1600 175
1600 8
926 8
926 156
8 0 25 0 0 0 0 142 0 0 402 5
1633 184
1591 184
1591 18
941 18
941 174
2 0 130 0 0 4224 0 128 0 0 273 3
1588 57
1625 57
1625 87
0 17 130 0 0 0 0 0 142 0 0 3
1625 84
1625 112
1627 112
1 17 131 0 0 8192 0 128 141 0 0 4
1552 57
1549 57
1549 330
1614 330
13 0 132 0 0 8320 0 142 0 0 279 3
1697 157
1700 157
1700 271
14 0 133 0 0 8192 0 142 0 0 280 4
1697 166
1718 166
1718 256
1723 256
15 0 134 0 0 8192 0 142 0 0 281 4
1697 175
1737 175
1737 243
1742 243
16 0 135 0 0 4096 0 142 0 0 282 4
1697 184
1759 184
1759 233
1764 233
13 4 132 0 0 0 0 141 140 0 0 4
1684 375
1700 375
1700 267
1772 267
14 3 133 0 0 8320 0 141 140 0 0 4
1684 384
1723 384
1723 255
1772 255
15 2 134 0 0 8320 0 141 140 0 0 4
1684 393
1742 393
1742 243
1772 243
16 1 135 0 0 8320 0 141 140 0 0 4
1684 402
1764 402
1764 231
1772 231
11 5 136 0 0 12416 0 135 141 0 0 4
1535 388
1542 388
1542 375
1620 375
9 6 137 0 0 12416 0 135 141 0 0 4
1535 352
1554 352
1554 384
1620 384
11 7 138 0 0 8320 0 134 141 0 0 4
1534 179
1564 179
1564 393
1620 393
9 8 139 0 0 8320 0 134 141 0 0 4
1534 143
1578 143
1578 402
1620 402
0 9 48 0 0 0 0 0 140 333 0 5
1219 924
1506 924
1506 486
1796 486
1796 297
8 1 7 0 0 0 0 140 139 0 0 3
1820 267
1917 267
1917 213
7 1 8 0 0 0 0 140 138 0 0 3
1820 255
1892 255
1892 213
6 1 9 0 0 0 0 140 137 0 0 3
1820 243
1863 243
1863 213
5 1 10 0 0 0 0 140 136 0 0 3
1820 231
1835 231
1835 213
1 3 127 0 0 4224 0 131 135 0 0 3
1316 364
1465 364
1465 361
8 0 125 0 0 0 0 135 0 0 305 4
1465 406
1394 406
1394 404
1396 404
7 1 126 0 0 12416 0 135 132 0 0 5
1465 397
1433 397
1433 463
1319 463
1319 464
6 0 125 0 0 0 0 135 0 0 305 2
1471 388
1396 388
5 0 125 0 0 0 0 135 0 0 305 2
1471 379
1396 379
4 0 125 0 0 0 0 135 0 0 305 4
1465 370
1401 370
1401 371
1396 371
2 0 125 0 0 0 0 135 0 0 305 2
1471 352
1396 352
1 0 125 0 0 0 0 135 0 0 305 2
1471 343
1396 343
6 0 125 0 0 0 0 134 0 0 305 2
1470 179
1396 179
5 0 125 0 0 0 0 134 0 0 305 2
1470 170
1396 170
4 0 125 0 0 0 0 134 0 0 305 4
1464 161
1400 161
1400 162
1396 162
2 0 125 0 0 0 0 134 0 0 305 2
1470 143
1396 143
1 0 125 0 0 0 0 134 0 0 305 2
1470 134
1396 134
1 18 125 0 0 12416 0 129 141 0 0 7
1396 80
1396 79
1396 79
1396 449
1688 449
1688 330
1684 330
2 1 140 0 0 4224 0 143 148 0 0 4
293 1033
494 1033
494 1183
514 1183
0 1 141 0 0 4096 0 0 143 332 0 7
665 841
400 841
400 984
221 984
221 1032
257 1032
257 1033
2 0 142 0 0 12416 0 148 0 0 310 5
520 1192
444 1192
444 1050
245 1050
245 1140
2 0 2 0 0 0 0 208 0 0 349 2
293 1140
357 1140
1 1 142 0 0 0 0 144 208 0 0 3
230 1139
230 1140
257 1140
2 0 143 0 0 4096 0 144 0 0 352 2
196 1139
163 1139
1 0 22 0 0 0 0 145 0 0 315 2
813 1295
813 1296
1 0 131 0 0 0 0 146 0 0 316 2
812 1208
812 1210
1 0 144 0 0 4096 0 147 0 0 317 2
815 1111
815 1114
4 0 22 0 0 24704 0 148 0 0 0 11
584 1219
676 1219
676 1296
1140 1296
1140 1373
316 1373
316 3221
538 3221
538 3170
549 3170
549 2420
5 1 131 0 0 16512 0 148 128 0 0 6
584 1210
1144 1210
1144 1177
1177 1177
1177 57
1552 57
6 0 144 0 0 12416 0 148 0 0 0 4
584 1201
677 1201
677 1114
1142 1114
7 3 145 0 0 12416 0 148 148 0 0 6
584 1192
627 1192
627 1082
470 1082
470 1210
520 1210
0 0 146 0 0 4096 0 0 0 378 336 2
721 475
721 915
2 2 147 0 0 4224 0 149 176 0 0 2
299 475
402 475
0 3 148 0 0 8320 0 0 176 380 0 5
824 457
824 619
350 619
350 493
402 493
0 1 149 0 0 12416 0 0 151 325 0 5
256 880
256 851
107 851
107 527
214 527
2 0 143 0 0 4096 0 150 0 0 352 2
212 879
163 879
2 0 2 0 0 0 0 209 0 0 349 4
300 879
353 879
353 881
358 881
1 1 149 0 0 0 0 150 209 0 0 5
246 879
246 880
256 880
256 879
264 879
2 1 150 0 0 12416 0 151 152 0 0 6
250 527
265 527
265 547
208 547
208 558
216 558
3 2 151 0 0 8320 0 152 164 0 0 6
261 567
326 567
326 392
260 392
260 352
287 352
0 2 13 0 0 12288 0 0 152 330 0 6
616 799
481 799
481 625
211 625
211 576
216 576
1 0 13 0 0 0 0 153 0 0 330 2
815 1050
815 1050
0 0 13 0 0 16512 0 0 0 379 12 9
767 466
767 799
611 799
611 1050
1538 1050
1538 1179
2414 1179
2414 1319
2711 1319
1 0 141 0 0 0 0 154 0 0 332 4
817 975
817 976
813 976
813 977
0 0 141 0 0 8192 0 0 0 354 0 3
665 709
665 977
1140 977
0 0 48 0 0 0 0 0 0 334 0 2
816 924
1227 924
1 3 48 0 0 0 0 155 156 0 0 3
816 922
816 924
792 924
2 0 152 0 0 4224 0 156 0 0 390 2
747 933
91 933
1 0 146 0 0 0 0 156 0 0 0 2
747 915
709 915
0 2 146 0 0 0 0 0 159 319 0 5
721 879
435 879
435 655
200 655
200 436
1 0 153 0 0 8320 0 158 0 0 340 5
187 386
130 386
130 820
255 820
255 841
2 0 2 0 0 0 0 210 0 0 349 2
298 841
358 841
1 1 153 0 0 0 0 157 210 0 0 3
246 842
246 841
262 841
2 0 143 0 0 0 0 157 0 0 352 2
212 842
163 842
3 3 154 0 0 8320 0 159 164 0 0 4
245 427
283 427
283 361
286 361
2 1 155 0 0 12416 0 158 159 0 0 6
223 386
250 386
250 401
193 401
193 418
200 418
1 3 156 0 0 4224 0 164 165 0 0 4
286 343
254 343
254 350
241 350
1 0 152 0 0 0 0 149 0 0 390 2
263 475
91 475
2 1 157 0 0 8320 0 160 165 0 0 5
211 297
211 315
179 315
179 341
196 341
0 1 158 0 0 12416 0 0 160 350 0 5
251 803
251 729
120 729
120 297
175 297
2 0 2 0 0 0 0 211 0 0 349 2
293 803
358 803
1 0 2 0 0 4224 0 161 0 0 0 4
357 1478
357 881
358 881
358 749
1 1 158 0 0 0 0 163 211 0 0 3
244 802
244 803
257 803
2 0 143 0 0 0 0 163 0 0 352 2
210 802
163 802
1 0 143 0 0 4224 0 162 0 0 0 2
163 770
163 1469
4 1 159 0 0 8320 0 164 176 0 0 4
332 352
391 352
391 466
396 466
2 0 141 0 0 12416 0 165 0 0 377 5
196 359
177 359
177 709
665 709
665 484
1 0 2 0 0 0 0 166 0 0 374 2
864 594
864 570
2 0 2 0 0 0 0 167 0 0 357 4
949 555
949 560
899 560
899 565
2 0 2 0 0 0 0 168 0 0 374 4
908 550
908 565
887 565
887 570
2 0 2 0 0 0 0 169 0 0 374 2
856 549
856 570
1 0 160 0 0 4096 0 167 0 0 383 4
949 535
949 435
922 435
922 430
1 0 161 0 0 4096 0 168 0 0 382 2
908 530
908 439
1 0 162 0 0 4096 0 169 0 0 381 2
856 529
856 448
1 0 148 0 0 0 0 170 0 0 380 2
802 531
802 457
1 0 13 0 0 0 0 171 0 0 379 2
744 525
744 466
1 0 146 0 0 0 0 172 0 0 378 2
685 525
685 475
1 0 141 0 0 0 0 173 0 0 377 2
625 524
625 484
1 0 163 0 0 4096 0 174 0 0 376 2
568 522
568 493
1 0 164 0 0 4096 0 175 0 0 375 2
509 521
509 502
2 0 2 0 0 0 0 170 0 0 374 2
802 551
802 570
2 0 2 0 0 0 0 171 0 0 374 2
744 545
744 570
2 0 2 0 0 0 0 172 0 0 374 2
685 545
685 570
2 0 2 0 0 0 0 173 0 0 374 2
625 544
625 570
2 0 2 0 0 0 0 174 0 0 374 2
568 542
568 570
2 0 2 0 0 0 0 175 0 0 374 2
509 541
509 570
0 0 2 0 0 0 0 0 0 0 0 2
482 570
894 570
4 0 164 0 0 4224 0 176 0 0 0 2
466 502
946 502
5 0 163 0 0 4096 0 176 0 0 0 2
466 493
959 493
6 0 141 0 0 0 0 176 0 0 0 2
466 484
947 484
7 0 146 0 0 4224 0 176 0 0 0 2
466 475
940 475
8 0 13 0 0 0 0 176 0 0 0 2
466 466
945 466
9 0 148 0 0 0 0 176 0 0 0 2
466 457
935 457
10 0 162 0 0 4224 0 176 0 0 0 2
466 448
940 448
11 0 161 0 0 4224 0 176 0 0 0 2
466 439
934 439
12 0 160 0 0 4224 0 176 0 0 0 2
466 430
929 430
13 0 165 0 0 4224 0 176 0 0 0 3
466 421
926 421
926 424
2 0 2 0 0 0 0 180 0 0 389 2
895 241
895 265
2 0 2 0 0 0 0 181 0 0 389 2
834 239
834 265
2 0 2 0 0 0 0 182 0 0 389 2
776 237
776 265
2 0 2 0 0 0 0 183 0 0 389 2
716 233
716 265
1 0 2 0 0 0 0 177 0 0 0 2
940 265
692 265
0 0 152 0 0 0 0 0 0 392 0 2
91 457
91 987
3 0 152 0 0 0 0 187 0 0 392 2
345 68
91 68
3 0 152 0 0 0 0 178 0 0 0 4
64 26
91 26
91 459
107 459
6 0 166 0 0 4096 0 184 0 0 394 2
620 174
527 174
11 0 166 0 0 4224 0 187 0 0 0 3
409 95
527 95
527 199
2 0 163 0 0 16512 0 179 0 0 376 7
168 172
158 172
158 171
150 171
150 680
587 680
587 493
1 0 152 0 0 0 0 179 0 0 392 5
168 154
168 127
237 127
237 80
91 80
2 3 167 0 0 12416 0 184 179 0 0 6
620 129
555 129
555 258
235 258
235 163
213 163
1 0 25 0 0 0 0 180 0 0 402 2
895 221
895 174
1 0 26 0 0 0 0 181 0 0 403 2
834 219
834 156
1 0 104 0 0 0 0 182 0 0 404 2
776 217
776 138
1 0 105 0 0 0 0 183 0 0 405 2
716 213
716 120
13 0 25 0 0 0 0 184 0 0 0 2
684 174
999 174
11 0 26 0 0 0 0 184 0 0 0 2
684 156
989 156
9 0 104 0 0 0 0 184 0 0 0 2
684 138
1130 138
7 0 105 0 0 0 0 184 0 0 0 2
684 120
1131 120
5 0 168 0 0 4224 0 184 0 0 414 2
620 165
479 165
4 0 169 0 0 4224 0 184 0 0 415 2
620 156
413 156
3 0 170 0 0 4224 0 184 0 0 416 2
620 147
355 147
1 0 171 0 0 12288 0 184 0 0 413 6
614 120
597 120
597 55
507 55
507 50
495 50
1 0 171 0 0 0 0 187 0 0 411 3
345 50
330 50
330 7
2 0 171 0 0 12416 0 187 0 0 413 5
345 59
309 59
309 7
461 7
461 50
9 0 171 0 0 0 0 187 0 0 413 3
415 59
489 59
489 50
8 1 171 0 0 0 0 187 185 0 0 4
415 50
495 50
495 39
503 39
0 12 168 0 0 0 0 0 187 0 0 3
479 172
479 104
409 104
0 13 169 0 0 0 0 0 187 0 0 5
413 172
413 141
428 141
428 113
409 113
0 14 170 0 0 0 0 0 187 0 0 5
355 169
355 136
423 136
423 122
409 122
0 1 2 0 0 0 0 0 186 418 0 5
345 118
262 118
262 175
268 175
268 188
7 6 2 0 0 0 0 187 187 0 0 2
345 122
345 113
5 6 2 0 0 0 0 187 187 0 0 2
345 104
345 113
4 5 2 0 0 0 0 187 187 0 0 2
345 95
345 104
21
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2786 1405 2863 1429
2797 1413 2851 1429
9 CORRECT !
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
2792 1573 2857 1597
2803 1581 2845 1597
7 WRONG !
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
2691 1257 2798 1281
2702 1264 2786 1280
14 Output Enabled
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2177 1254 2202 1278
2185 1262 2193 1278
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1971 1257 1996 1281
1979 1265 1987 1281
1 N
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1926 1233 2043 1257
1936 1241 2032 1257
12 FIRST NUMBER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
2137 1232 2262 1256
2147 1240 2251 1256
13 SECOND NUMBER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
435 818 649 841
447 828 636 843
27 Question Mode Change Enable
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 38
1155 1275 1448 1298
1168 1285 1434 1300
38 To master/slave selector of Expression
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
1148 1191 1455 1214
1161 1201 1441 1216
40 To master/slave selector of Venn Diagram
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
901 1269 1061 1292
914 1279 1047 1294
19 Expression Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
900 1182 1073 1205
912 1192 1060 1207
21 Venn Diagram Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
901 1084 984 1107
914 1094 970 1109
8 DIY Mode
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
477 655 630 678
490 665 616 680
18 Load Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
-11 68 100 91
2 78 86 93
12 Clock Signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
457 327 603 350
470 337 589 352
17 Master Controller
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
870 1016 1035 1039
882 1026 1022 1041
20 Output Enable signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
871 86 987 109
883 96 974 111
13 Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
610 10 796 33
622 20 783 35
23 Random Number Generator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
871 948 1050 971
883 958 1037 973
22 Reset signal for slave
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
870 893 1049 916
882 903 1036 918
22 Master Clock for Slave
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
