CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 60 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
37 D:\Programs\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.209790 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
69
7 Ground~
168 1209 520 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
5.90066e-315 0
0
5 4049~
219 1567 57 0 2 22
0 13 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
391 0 0
2
5.90066e-315 0
0
2 +V
167 1396 71 0 1 3
0 3
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.90066e-315 0
0
14 NO PushButton~
191 1303 146 0 2 5
0 7 2
0
0 0 4720 0
0
2 S9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3421 0 0
2
5.90066e-315 5.42933e-315
0
14 NO PushButton~
191 1299 356 0 2 5
0 5 2
0
0 0 4720 0
0
2 S8
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8157 0 0
2
5.90066e-315 5.41896e-315
0
14 NO PushButton~
191 1302 456 0 2 5
0 4 2
0
0 0 4720 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5572 0 0
2
5.90066e-315 5.41378e-315
0
14 NO PushButton~
191 1300 251 0 2 5
0 6 2
0
0 0 4720 0
0
2 S6
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8901 0 0
2
5.90066e-315 5.4086e-315
0
6 74LS73
102 1502 161 0 12 25
0 3 3 7 3 3 3 6 3 21
61 20 62
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
3 U15
-10 -52 11 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
5.90066e-315 5.40342e-315
0
6 74LS73
102 1503 370 0 12 25
0 3 3 5 3 3 3 4 3 19
63 18 64
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
3 U14
-10 -52 11 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.90066e-315 5.39824e-315
0
14 Logic Display~
6 1835 195 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90066e-315 5.39306e-315
0
14 Logic Display~
6 1863 195 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90066e-315 5.38788e-315
0
14 Logic Display~
6 1892 195 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.90066e-315 5.37752e-315
0
14 Logic Display~
6 1917 195 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.90066e-315 5.36716e-315
0
12 Quad D Flop~
47 1796 261 0 9 19
0 17 16 15 14 26 25 24 23 22
0
0 0 4720 0
4 QDFF
-14 -44 14 -36
3 U13
-10 -46 11 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4597 0 0
2
5.90066e-315 5.3568e-315
0
7 74LS245
64 1652 366 0 18 37
0 65 66 67 68 18 19 20 21 69
70 71 72 14 15 16 17 13 3
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
3 U12
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
3835 0 0
2
5.90066e-315 5.32571e-315
0
7 74LS245
64 1665 148 0 18 37
0 73 74 75 76 8 9 10 11 77
78 79 80 14 15 16 17 12 3
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
3 U11
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
5.90066e-315 5.30499e-315
0
5 4049~
219 272 1033 0 2 22
0 28 27
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
5616 0 0
2
44974.8 0
0
14 NO PushButton~
191 213 1131 0 2 5
0 29 30
0
0 0 4720 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9323 0 0
2
44974.8 1
0
14 Logic Display~
6 813 1277 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
44974.8 2
0
14 Logic Display~
6 812 1190 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44974.8 3
0
14 Logic Display~
6 815 1093 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
44974.8 4
0
4 4017
219 552 1165 0 14 29
0 27 29 33 31 13 32 33 81 82
83 84 85 86 87
0
0 0 6896 0
4 4017
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
9672 0 0
2
44974.8 5
0
5 4049~
219 278 475 0 2 22
0 41 35
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
7876 0 0
2
44974.8 6
0
14 NO PushButton~
191 229 871 0 2 5
0 37 30
0
0 0 4720 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6369 0 0
2
44974.8 7
0
5 4049~
219 229 527 0 2 22
0 37 38
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
9172 0 0
2
44974.8 8
0
9 2-In AND~
219 240 567 0 3 22
0 38 40 39
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7100 0 0
2
44974.8 9
0
14 Logic Display~
6 815 1032 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
44974.8 10
0
14 Logic Display~
6 817 957 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
44974.8 11
0
14 Logic Display~
6 816 904 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90066e-315 0
0
9 2-In AND~
219 771 924 0 3 22
0 34 41 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3178 0 0
2
5.90066e-315 5.26354e-315
0
14 NO PushButton~
191 229 834 0 2 5
0 42 30
0
0 0 4720 0
0
2 S2
-7 -22 7 -14
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3409 0 0
2
5.90066e-315 5.30499e-315
0
5 4049~
219 202 386 0 2 22
0 42 44
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
3951 0 0
2
5.90066e-315 5.32571e-315
0
9 2-In AND~
219 224 427 0 3 22
0 44 34 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8885 0 0
2
5.90066e-315 5.34643e-315
0
5 4049~
219 190 297 0 2 22
0 47 46
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3780 0 0
2
5.90066e-315 5.3568e-315
0
7 Ground~
168 357 1484 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
5.90066e-315 5.36716e-315
0
2 +V
167 163 761 0 1 3
0 30
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
5.90066e-315 5.37752e-315
0
14 NO PushButton~
191 227 794 0 2 5
0 47 30
0
0 0 4720 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9424 0 0
2
5.90066e-315 5.38788e-315
0
8 3-In OR~
219 299 352 0 4 22
0 45 39 43 48
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
9968 0 0
2
5.90066e-315 5.39306e-315
0
9 2-In AND~
219 220 350 0 3 22
0 46 28 45
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9281 0 0
2
5.90066e-315 5.39824e-315
0
7 Ground~
168 864 600 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8464 0 0
2
5.90066e-315 5.40342e-315
0
4 LED~
171 949 545 0 2 2
10 49 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D13
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7168 0 0
2
5.90066e-315 5.4086e-315
0
4 LED~
171 908 540 0 2 2
10 50 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D12
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3171 0 0
2
5.90066e-315 5.41378e-315
0
4 LED~
171 856 539 0 2 2
10 51 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D11
20 -10 41 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4139 0 0
2
5.90066e-315 5.41896e-315
0
4 LED~
171 802 541 0 2 2
10 36 2
0
0 0 880 0
4 LED1
17 0 45 8
3 D10
21 -10 42 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6435 0 0
2
5.90066e-315 5.42414e-315
0
4 LED~
171 744 535 0 2 2
10 40 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D9
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5283 0 0
2
5.90066e-315 5.42933e-315
0
4 LED~
171 685 535 0 2 2
10 34 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6874 0 0
2
5.90066e-315 5.43192e-315
0
4 LED~
171 625 534 0 2 2
10 28 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5305 0 0
2
5.90066e-315 5.43451e-315
0
4 LED~
171 568 532 0 2 2
10 52 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
34 0 0
2
5.90066e-315 5.4371e-315
0
4 LED~
171 509 531 0 2 2
10 53 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
969 0 0
2
5.90066e-315 5.43969e-315
0
4 4017
219 434 448 0 14 29
0 48 35 36 53 52 28 34 40 36
51 50 49 54 88
0
0 0 6896 0
4 4017
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
102 %D [%16bi %8bi %1i %2i %3i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 13 14 15 3 2 4 7 10 1
5 6 9 11 12 13 14 15 3 2
4 7 10 1 5 6 9 11 12 0
65 0 0 512 1 0 0 0
1 U
8402 0 0
2
5.90066e-315 5.44228e-315
0
7 Ground~
168 940 271 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3751 0 0
2
5.90066e-315 5.44487e-315
0
7 Pulser~
4 40 35 0 10 12
0 89 90 41 91 0 0 5 5 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4292 0 0
2
5.90066e-315 5.44746e-315
0
9 2-In AND~
219 192 163 0 3 22
0 41 52 56
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6118 0 0
2
44974.8 12
0
4 LED~
171 895 231 0 2 2
10 11 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
34 0 0
2
44974.8 13
0
4 LED~
171 834 229 0 2 2
10 10 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6357 0 0
2
44974.8 14
0
4 LED~
171 776 227 0 2 2
10 9 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
319 0 0
2
44974.8 15
0
4 LED~
171 716 223 0 2 2
10 8 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3976 0 0
2
44974.8 16
0
7 74LS175
131 652 147 0 14 29
0 60 56 59 58 57 55 8 92 9
93 10 94 11 95
0
0 0 4848 0
7 74LS175
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 9 13 12 5 4 15 14 10
11 7 6 2 3 1 9 13 12 5
4 15 14 10 11 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
7634 0 0
2
44974.8 17
0
2 +V
167 503 30 0 1 3
0 60
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
523 0 0
2
44974.8 18
0
7 Ground~
168 268 194 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6748 0 0
2
44974.8 19
0
7 74LS161
96 377 86 0 14 29
0 60 60 41 2 2 2 2 60 60
96 55 57 58 59
0
0 0 6896 0
8 74LS161A
-28 -60 28 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
6901 0 0
2
44974.8 20
0
9 Resistor~
219 1355 440 0 4 5
0 4 3 0 1
0
0 0 880 0
2 1k
-7 -15 7 -7
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
842 0 0
2
5.90066e-315 0
0
9 Resistor~
219 1348 336 0 4 5
0 5 3 0 1
0
0 0 880 0
2 1k
-7 -15 7 -7
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3277 0 0
2
5.90066e-315 0
0
9 Resistor~
219 1335 220 0 4 5
0 6 3 0 1
0
0 0 880 0
2 1k
-7 -15 7 -7
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4212 0 0
2
5.90066e-315 0
0
9 Resistor~
219 1347 117 0 4 5
0 7 3 0 1
0
0 0 880 0
2 1k
-7 -15 7 -7
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4720 0 0
2
5.90066e-315 0
0
9 Resistor~
219 275 1140 0 4 5
0 29 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5551 0 0
2
44974.8 21
0
9 Resistor~
219 282 879 0 4 5
0 37 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R4
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6986 0 0
2
44974.8 22
0
9 Resistor~
219 280 841 0 4 5
0 42 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-8 -26 6 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8745 0 0
2
5.90066e-315 5.45005e-315
0
9 Resistor~
219 275 803 0 4 5
0 47 2 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-9 -24 5 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9592 0 0
2
44974.8 23
0
171
0 18 3 0 0 4096 0 0 16 55 0 4
1396 244
1731 244
1731 112
1697 112
2 0 3 0 0 0 0 62 0 0 55 2
1373 440
1396 440
2 0 3 0 0 0 0 63 0 0 55 2
1366 336
1396 336
2 0 3 0 0 0 0 64 0 0 55 2
1353 220
1396 220
2 0 3 0 0 0 0 65 0 0 55 2
1365 117
1396 117
1 0 4 0 0 4096 0 62 0 0 44 2
1337 440
1337 463
1 0 5 0 0 4096 0 63 0 0 42 2
1330 336
1330 364
1 1 6 0 0 4096 0 64 7 0 0 2
1317 220
1317 259
1 0 7 0 0 4096 0 65 0 0 14 2
1329 117
1329 152
2 0 2 0 0 4096 0 6 0 0 16 2
1285 464
1209 464
2 0 2 0 0 0 0 5 0 0 16 2
1282 364
1209 364
1 7 6 0 0 12416 0 7 8 0 0 4
1317 259
1363 259
1363 188
1464 188
2 0 2 0 0 0 0 7 0 0 16 2
1283 259
1209 259
1 3 7 0 0 8320 0 4 8 0 0 3
1320 154
1320 152
1464 152
2 0 2 0 0 4096 0 4 0 0 16 2
1286 154
1209 154
0 1 2 0 0 4096 0 0 1 0 0 2
1209 71
1209 514
8 0 3 0 0 0 0 8 0 0 55 2
1464 197
1396 197
5 0 8 0 0 12416 0 16 0 0 156 5
1633 157
1614 157
1614 41
893 41
893 120
6 0 9 0 0 12416 0 16 0 0 155 5
1633 166
1608 166
1608 30
912 30
912 138
7 0 10 0 0 12416 0 16 0 0 154 5
1633 175
1600 175
1600 8
926 8
926 156
8 0 11 0 0 12416 0 16 0 0 153 5
1633 184
1591 184
1591 18
941 18
941 174
2 0 12 0 0 4224 0 2 0 0 23 3
1588 57
1625 57
1625 87
0 17 12 0 0 0 0 0 16 0 0 3
1625 84
1625 112
1627 112
1 17 13 0 0 8192 0 2 15 0 0 4
1552 57
1549 57
1549 330
1614 330
13 0 14 0 0 8320 0 16 0 0 29 3
1697 157
1700 157
1700 271
14 0 15 0 0 8192 0 16 0 0 30 4
1697 166
1718 166
1718 256
1723 256
15 0 16 0 0 8192 0 16 0 0 31 4
1697 175
1737 175
1737 243
1742 243
16 0 17 0 0 4096 0 16 0 0 32 4
1697 184
1759 184
1759 233
1764 233
13 4 14 0 0 0 0 15 14 0 0 4
1684 375
1700 375
1700 267
1772 267
14 3 15 0 0 8320 0 15 14 0 0 4
1684 384
1723 384
1723 255
1772 255
15 2 16 0 0 8320 0 15 14 0 0 4
1684 393
1742 393
1742 243
1772 243
16 1 17 0 0 8320 0 15 14 0 0 4
1684 402
1764 402
1764 231
1772 231
11 5 18 0 0 12416 0 9 15 0 0 4
1535 388
1542 388
1542 375
1620 375
9 6 19 0 0 12416 0 9 15 0 0 4
1535 352
1554 352
1554 384
1620 384
11 7 20 0 0 8320 0 8 15 0 0 4
1534 179
1564 179
1564 393
1620 393
9 8 21 0 0 8320 0 8 15 0 0 4
1534 143
1578 143
1578 402
1620 402
0 9 22 0 0 8320 0 0 14 84 0 5
1219 924
1506 924
1506 486
1796 486
1796 297
8 1 23 0 0 4224 0 14 13 0 0 3
1820 267
1917 267
1917 213
7 1 24 0 0 4224 0 14 12 0 0 3
1820 255
1892 255
1892 213
6 1 25 0 0 4224 0 14 11 0 0 3
1820 243
1863 243
1863 213
5 1 26 0 0 8320 0 14 10 0 0 3
1820 231
1835 231
1835 213
1 3 5 0 0 4224 0 5 9 0 0 3
1316 364
1465 364
1465 361
8 0 3 0 0 0 0 9 0 0 55 4
1465 406
1394 406
1394 404
1396 404
7 1 4 0 0 12416 0 9 6 0 0 5
1465 397
1433 397
1433 463
1319 463
1319 464
6 0 3 0 0 0 0 9 0 0 55 2
1471 388
1396 388
5 0 3 0 0 0 0 9 0 0 55 2
1471 379
1396 379
4 0 3 0 0 0 0 9 0 0 55 4
1465 370
1401 370
1401 371
1396 371
2 0 3 0 0 0 0 9 0 0 55 2
1471 352
1396 352
1 0 3 0 0 0 0 9 0 0 55 2
1471 343
1396 343
6 0 3 0 0 0 0 8 0 0 55 2
1470 179
1396 179
5 0 3 0 0 0 0 8 0 0 55 2
1470 170
1396 170
4 0 3 0 0 0 0 8 0 0 55 4
1464 161
1400 161
1400 162
1396 162
2 0 3 0 0 0 0 8 0 0 55 2
1470 143
1396 143
1 0 3 0 0 0 0 8 0 0 55 2
1470 134
1396 134
1 18 3 0 0 12416 0 3 15 0 0 7
1396 80
1396 79
1396 79
1396 449
1688 449
1688 330
1684 330
0 0 2 0 0 4224 0 0 0 0 100 4
1227 887
466 887
466 1014
357 1014
2 1 27 0 0 4224 0 17 22 0 0 4
293 1033
494 1033
494 1183
514 1183
0 1 28 0 0 4096 0 0 17 83 0 7
665 841
400 841
400 984
221 984
221 1032
257 1032
257 1033
2 0 29 0 0 12416 0 22 0 0 61 5
520 1192
444 1192
444 1050
245 1050
245 1140
2 0 2 0 0 0 0 66 0 0 100 2
293 1140
357 1140
1 1 29 0 0 0 0 18 66 0 0 3
230 1139
230 1140
257 1140
2 0 30 0 0 4096 0 18 0 0 103 2
196 1139
163 1139
1 0 31 0 0 4096 0 19 0 0 66 2
813 1295
813 1296
1 0 13 0 0 0 0 20 0 0 67 2
812 1208
812 1210
1 0 32 0 0 4096 0 21 0 0 68 2
815 1111
815 1114
4 0 31 0 0 12416 0 22 0 0 0 4
584 1219
676 1219
676 1296
1142 1296
5 1 13 0 0 16512 0 22 2 0 0 6
584 1210
1144 1210
1144 1177
1177 1177
1177 57
1552 57
6 0 32 0 0 12416 0 22 0 0 0 4
584 1201
677 1201
677 1114
1142 1114
7 3 33 0 0 12416 0 22 22 0 0 6
584 1192
627 1192
627 1082
470 1082
470 1210
520 1210
0 0 34 0 0 4096 0 0 0 129 87 2
721 475
721 915
2 2 35 0 0 4224 0 23 50 0 0 2
299 475
402 475
0 3 36 0 0 8320 0 0 50 131 0 5
824 457
824 619
350 619
350 493
402 493
0 1 37 0 0 12416 0 0 25 76 0 5
256 880
256 851
107 851
107 527
214 527
2 0 30 0 0 4096 0 24 0 0 103 2
212 879
163 879
2 0 2 0 0 0 0 67 0 0 100 4
300 879
353 879
353 881
358 881
1 1 37 0 0 0 0 24 67 0 0 5
246 879
246 880
256 880
256 879
264 879
2 1 38 0 0 12416 0 25 26 0 0 6
250 527
265 527
265 547
208 547
208 558
216 558
3 2 39 0 0 8320 0 26 38 0 0 6
261 567
326 567
326 392
260 392
260 352
287 352
0 2 40 0 0 12288 0 0 26 81 0 6
616 799
481 799
481 625
211 625
211 576
216 576
1 0 40 0 0 0 0 27 0 0 81 2
815 1050
815 1050
0 0 40 0 0 16512 0 0 0 130 0 5
767 466
767 799
611 799
611 1050
1141 1050
1 0 28 0 0 0 0 28 0 0 83 4
817 975
817 976
813 976
813 977
0 0 28 0 0 8192 0 0 0 105 0 3
665 709
665 977
1140 977
0 0 22 0 0 0 0 0 0 85 0 2
816 924
1227 924
1 3 22 0 0 0 0 29 30 0 0 3
816 922
816 924
792 924
2 0 41 0 0 4224 0 30 0 0 141 2
747 933
91 933
1 0 34 0 0 0 0 30 0 0 0 2
747 915
709 915
0 2 34 0 0 0 0 0 33 70 0 5
721 879
435 879
435 655
200 655
200 436
1 0 42 0 0 8320 0 32 0 0 91 5
187 386
130 386
130 820
255 820
255 841
2 0 2 0 0 0 0 68 0 0 100 2
298 841
358 841
1 1 42 0 0 0 0 31 68 0 0 3
246 842
246 841
262 841
2 0 30 0 0 0 0 31 0 0 103 2
212 842
163 842
3 3 43 0 0 8320 0 33 38 0 0 4
245 427
283 427
283 361
286 361
2 1 44 0 0 12416 0 32 33 0 0 6
223 386
250 386
250 401
193 401
193 418
200 418
1 3 45 0 0 4224 0 38 39 0 0 4
286 343
254 343
254 350
241 350
1 0 41 0 0 0 0 23 0 0 141 2
263 475
91 475
2 1 46 0 0 8320 0 34 39 0 0 5
211 297
211 315
179 315
179 341
196 341
0 1 47 0 0 12416 0 0 34 101 0 5
251 803
251 729
120 729
120 297
175 297
2 0 2 0 0 0 0 69 0 0 100 2
293 803
358 803
1 0 2 0 0 0 0 35 0 0 0 4
357 1478
357 881
358 881
358 749
1 1 47 0 0 0 0 37 69 0 0 3
244 802
244 803
257 803
2 0 30 0 0 0 0 37 0 0 103 2
210 802
163 802
1 0 30 0 0 4224 0 36 0 0 0 2
163 770
163 1469
4 1 48 0 0 8320 0 38 50 0 0 4
332 352
391 352
391 466
396 466
2 0 28 0 0 12416 0 39 0 0 128 5
196 359
177 359
177 709
665 709
665 484
1 0 2 0 0 0 0 40 0 0 125 2
864 594
864 570
2 0 2 0 0 0 0 41 0 0 108 4
949 555
949 560
899 560
899 565
2 0 2 0 0 0 0 42 0 0 125 4
908 550
908 565
887 565
887 570
2 0 2 0 0 0 0 43 0 0 125 2
856 549
856 570
1 0 49 0 0 4096 0 41 0 0 134 4
949 535
949 435
922 435
922 430
1 0 50 0 0 4096 0 42 0 0 133 2
908 530
908 439
1 0 51 0 0 4096 0 43 0 0 132 2
856 529
856 448
1 0 36 0 0 0 0 44 0 0 131 2
802 531
802 457
1 0 40 0 0 0 0 45 0 0 130 2
744 525
744 466
1 0 34 0 0 0 0 46 0 0 129 2
685 525
685 475
1 0 28 0 0 0 0 47 0 0 128 2
625 524
625 484
1 0 52 0 0 4096 0 48 0 0 127 2
568 522
568 493
1 0 53 0 0 4096 0 49 0 0 126 2
509 521
509 502
2 0 2 0 0 0 0 44 0 0 125 2
802 551
802 570
2 0 2 0 0 0 0 45 0 0 125 2
744 545
744 570
2 0 2 0 0 0 0 46 0 0 125 2
685 545
685 570
2 0 2 0 0 0 0 47 0 0 125 2
625 544
625 570
2 0 2 0 0 0 0 48 0 0 125 2
568 542
568 570
2 0 2 0 0 0 0 49 0 0 125 2
509 541
509 570
0 0 2 0 0 0 0 0 0 0 0 2
482 570
894 570
4 0 53 0 0 4224 0 50 0 0 0 2
466 502
946 502
5 0 52 0 0 4096 0 50 0 0 0 2
466 493
959 493
6 0 28 0 0 0 0 50 0 0 0 2
466 484
947 484
7 0 34 0 0 4224 0 50 0 0 0 2
466 475
940 475
8 0 40 0 0 0 0 50 0 0 0 2
466 466
945 466
9 0 36 0 0 0 0 50 0 0 0 2
466 457
935 457
10 0 51 0 0 4224 0 50 0 0 0 2
466 448
940 448
11 0 50 0 0 4224 0 50 0 0 0 2
466 439
934 439
12 0 49 0 0 4224 0 50 0 0 0 2
466 430
929 430
13 0 54 0 0 4224 0 50 0 0 0 3
466 421
926 421
926 424
2 0 2 0 0 0 0 54 0 0 140 2
895 241
895 265
2 0 2 0 0 0 0 55 0 0 140 2
834 239
834 265
2 0 2 0 0 0 0 56 0 0 140 2
776 237
776 265
2 0 2 0 0 0 0 57 0 0 140 2
716 233
716 265
1 0 2 0 0 0 0 51 0 0 0 2
940 265
692 265
0 0 41 0 0 0 0 0 0 143 0 2
91 457
91 987
3 0 41 0 0 0 0 61 0 0 143 2
345 68
91 68
3 0 41 0 0 0 0 52 0 0 0 4
64 26
91 26
91 459
107 459
6 0 55 0 0 4096 0 58 0 0 145 2
620 174
527 174
11 0 55 0 0 4224 0 61 0 0 0 3
409 95
527 95
527 199
2 0 52 0 0 16512 0 53 0 0 127 7
168 172
158 172
158 171
150 171
150 680
587 680
587 493
1 0 41 0 0 0 0 53 0 0 143 5
168 154
168 127
237 127
237 80
91 80
2 3 56 0 0 12416 0 58 53 0 0 6
620 129
555 129
555 258
235 258
235 163
213 163
1 0 11 0 0 0 0 54 0 0 153 2
895 221
895 174
1 0 10 0 0 0 0 55 0 0 154 2
834 219
834 156
1 0 9 0 0 0 0 56 0 0 155 2
776 217
776 138
1 0 8 0 0 0 0 57 0 0 156 2
716 213
716 120
13 0 11 0 0 0 0 58 0 0 0 2
684 174
999 174
11 0 10 0 0 0 0 58 0 0 0 2
684 156
989 156
9 0 9 0 0 0 0 58 0 0 0 2
684 138
975 138
7 0 8 0 0 0 0 58 0 0 0 2
684 120
961 120
5 0 57 0 0 4224 0 58 0 0 165 2
620 165
479 165
4 0 58 0 0 4224 0 58 0 0 166 2
620 156
413 156
3 0 59 0 0 4224 0 58 0 0 167 2
620 147
355 147
1 0 60 0 0 12288 0 58 0 0 164 6
614 120
597 120
597 55
507 55
507 50
495 50
1 0 60 0 0 0 0 61 0 0 162 3
345 50
330 50
330 7
2 0 60 0 0 12416 0 61 0 0 164 5
345 59
309 59
309 7
461 7
461 50
9 0 60 0 0 0 0 61 0 0 164 3
415 59
489 59
489 50
8 1 60 0 0 0 0 61 59 0 0 4
415 50
495 50
495 39
503 39
0 12 57 0 0 0 0 0 61 0 0 3
479 172
479 104
409 104
0 13 58 0 0 0 0 0 61 0 0 5
413 172
413 141
428 141
428 113
409 113
0 14 59 0 0 0 0 0 61 0 0 5
355 169
355 136
423 136
423 122
409 122
0 1 2 0 0 0 0 0 60 169 0 5
345 118
262 118
262 175
268 175
268 188
7 6 2 0 0 0 0 61 61 0 0 2
345 122
345 113
5 6 2 0 0 0 0 61 61 0 0 2
345 104
345 113
4 5 2 0 0 0 0 61 61 0 0 2
345 95
345 104
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
435 818 649 841
447 828 636 843
27 Question Mode Change Enable
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 38
1155 1275 1448 1298
1168 1285 1434 1300
38 To master/slave selector of Expression
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
1148 1191 1455 1214
1161 1201 1441 1216
40 To master/slave selector of Venn Diagram
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
901 1269 1061 1292
914 1279 1047 1294
19 Expression Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
900 1182 1073 1205
912 1192 1060 1207
21 Venn Diagram Question
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
901 1084 984 1107
914 1094 970 1109
8 DIY Mode
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
477 655 630 678
490 665 616 680
18 Load Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
-11 68 100 91
2 78 86 93
12 Clock Signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
457 327 603 350
470 337 589 352
17 Master Controller
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
870 1016 1035 1039
882 1026 1022 1041
20 Output Enable signal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
871 86 987 109
883 96 974 111
13 Random Number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
610 10 796 33
622 20 783 35
23 Random Number Generator
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
871 948 1050 971
883 958 1037 973
22 Reset signal for slave
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
870 893 1049 916
882 903 1036 918
22 Master Clock for Slave
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
