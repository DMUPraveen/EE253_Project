CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 50 10
78 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
246 176 359 273
9437202 0
0
6 Title:
5 Name:
0
0
0
128
13 Logic Switch~
5 787 1274 0 1 11
0 92
0
0 0 21344 90
2 0V
14 0 28 8
2 M0
14 -10 28 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9796 0 0
2
5.90066e-315 0
0
13 Logic Switch~
5 716 1272 0 1 11
0 93
0
0 0 21344 90
2 0V
14 0 28 8
2 M1
12 -13 26 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5952 0 0
2
5.90066e-315 5.26354e-315
0
13 Logic Switch~
5 653 1272 0 1 11
0 94
0
0 0 21344 90
2 0V
14 0 28 8
2 M2
13 -10 27 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3649 0 0
2
5.90066e-315 5.30499e-315
0
13 Logic Switch~
5 591 1275 0 1 11
0 95
0
0 0 21344 90
2 0V
14 0 28 8
2 M3
14 -10 28 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3716 0 0
2
5.90066e-315 5.32571e-315
0
13 Logic Switch~
5 528 1272 0 1 11
0 32
0
0 0 21344 90
2 0V
14 0 28 8
1 S
17 -10 24 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4797 0 0
2
5.90066e-315 5.34643e-315
0
13 Logic Switch~
5 1456 837 0 1 11
0 53
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4681 0 0
2
5.90066e-315 5.3568e-315
0
13 Logic Switch~
5 1456 874 0 1 11
0 52
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9730 0 0
2
5.90066e-315 5.36716e-315
0
2 +V
167 1822 78 0 1 3
0 7
0
0 0 54240 0
3 15V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9874 0 0
2
44974.8 0
0
14 NO PushButton~
191 1961 239 0 2 5
0 5 7
0
0 0 4704 0
0
3 S24
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
364 0 0
2
44974.8 1
0
14 NO PushButton~
191 1963 444 0 2 5
0 3 7
0
0 0 4704 0
0
3 S23
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3656 0 0
2
44974.8 2
0
14 NO PushButton~
191 1960 344 0 2 5
0 4 7
0
0 0 4704 0
0
3 S22
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3131 0 0
2
44974.8 3
0
7 Ground~
168 2007 555 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6772 0 0
2
44974.8 4
0
14 NO PushButton~
191 1964 134 0 2 5
0 6 7
0
0 0 4704 0
0
3 S21
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9557 0 0
2
44974.8 5
0
2 +V
167 1575 80 0 1 3
0 14
0
0 0 54240 0
3 15V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5789 0 0
2
44974.8 6
0
14 NO PushButton~
191 1714 241 0 2 5
0 12 14
0
0 0 4704 0
0
3 S20
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7328 0 0
2
44974.8 7
0
14 NO PushButton~
191 1716 446 0 2 5
0 10 14
0
0 0 4704 0
0
3 S19
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4799 0 0
2
44974.8 8
0
14 NO PushButton~
191 1713 346 0 2 5
0 11 14
0
0 0 4704 0
0
3 S18
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9196 0 0
2
44974.8 9
0
7 Ground~
168 1760 557 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3857 0 0
2
44974.8 10
0
14 NO PushButton~
191 1717 136 0 2 5
0 13 14
0
0 0 4704 0
0
3 S17
-11 -20 10 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7125 0 0
2
44974.8 11
0
14 NO PushButton~
191 165 810 0 2 5
0 20 21
0
0 0 4704 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3641 0 0
2
44974.8 12
0
7 Ground~
168 208 1231 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9821 0 0
2
44974.8 13
0
14 NO PushButton~
191 161 1020 0 2 5
0 18 21
0
0 0 4704 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3187 0 0
2
44974.8 14
0
14 NO PushButton~
191 164 1120 0 2 5
0 17 21
0
0 0 4704 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
762 0 0
2
44974.8 15
0
14 NO PushButton~
191 162 915 0 2 5
0 19 21
0
0 0 4704 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
39 0 0
2
44974.8 16
0
2 +V
167 33 66 0 1 3
0 21
0
0 0 54240 0
3 15V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9450 0 0
2
44974.8 17
0
14 NO PushButton~
191 172 227 0 2 5
0 24 21
0
0 0 4704 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3236 0 0
2
5.90066e-315 5.37752e-315
0
14 NO PushButton~
191 174 432 0 2 5
0 22 21
0
0 0 4704 0
0
2 S6
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3321 0 0
2
5.90066e-315 5.38788e-315
0
14 NO PushButton~
191 171 332 0 2 5
0 23 21
0
0 0 4704 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8879 0 0
2
5.90066e-315 5.39306e-315
0
7 Ground~
168 218 543 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5433 0 0
2
5.90066e-315 5.39824e-315
0
14 NO PushButton~
191 175 122 0 2 5
0 25 21
0
0 0 4704 0
0
2 S8
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3679 0 0
2
5.90066e-315 5.40342e-315
0
5 74148
219 694 388 0 14 29
0 2 36 37 38 39 40 41 42 43
2 35 34 33 27
0
0 0 6880 270
5 74148
-18 -60 17 -52
3 U10
56 -2 77 6
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 3 2 1 13 12 11 10
15 9 7 6 14 5 4 3 2 1
13 12 11 10 15 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
9342 0 0
2
5.90066e-315 5.4086e-315
0
7 74LS154
95 1578 929 0 22 45
0 53 52 89 88 87 86 54 55 56
57 58 59 60 61 62 63 64 65 66
67 68 69
0
0 0 4832 0
6 74F154
-21 -87 21 -79
2 U5
-7 -88 7 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
3623 0 0
2
5.90066e-315 5.41378e-315
0
9 Inverter~
13 662 493 0 2 22
0 35 31
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U3E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3722 0 0
2
5.90066e-315 5.41896e-315
0
9 Inverter~
13 693 494 0 2 22
0 34 91
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U3F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
8993 0 0
2
5.90066e-315 5.42414e-315
0
9 Inverter~
13 724 494 0 2 22
0 33 30
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3723 0 0
2
5.90066e-315 5.42933e-315
0
8 4-In OR~
219 1211 162 0 5 22
0 13 12 11 10 114
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
6244 0 0
2
5.90066e-315 5.43192e-315
0
8 4-In OR~
219 1213 241 0 5 22
0 6 5 4 3 113
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U4B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
6421 0 0
2
5.90066e-315 5.43451e-315
0
8 2-In OR~
219 1294 201 0 3 22
0 114 113 90
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7743 0 0
2
5.90066e-315 5.4371e-315
0
12 D Flip-Flop~
219 1186 1016 0 4 9
0 98 28 115 87
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U11
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9840 0 0
2
5.90066e-315 5.43969e-315
0
12 D Flip-Flop~
219 1188 1174 0 4 9
0 97 28 116 86
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U9
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6910 0 0
2
5.90066e-315 5.44228e-315
0
12 D Flip-Flop~
219 1183 849 0 4 9
0 99 28 117 88
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U8
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
449 0 0
2
5.90066e-315 5.44487e-315
0
12 D Flip-Flop~
219 1182 692 0 4 9
0 100 28 118 89
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8761 0 0
2
5.90066e-315 5.44746e-315
0
9 2-In AND~
219 975 664 0 3 22
0 90 95 111
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
6748 0 0
2
5.90066e-315 5.45005e-315
0
8 3-In OR~
219 1071 653 0 4 22
0 112 111 110 100
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 12 0
1 U
7393 0 0
2
5.90066e-315 5.45264e-315
0
9 2-In AND~
219 974 710 0 3 22
0 32 95 110
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
7699 0 0
2
5.90066e-315 5.45523e-315
0
9 2-In AND~
219 976 614 0 3 22
0 96 90 112
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
6638 0 0
2
5.90066e-315 5.45782e-315
0
9 2-In AND~
219 974 775 0 3 22
0 96 30 109
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
4595 0 0
2
5.90066e-315 5.46041e-315
0
9 2-In AND~
219 972 871 0 3 22
0 32 94 107
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U17A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
9395 0 0
2
5.90066e-315 5.463e-315
0
8 3-In OR~
219 1069 814 0 4 22
0 109 108 107 99
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U2B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 12 0
1 U
3303 0 0
2
5.90066e-315 5.46559e-315
0
9 2-In AND~
219 973 825 0 3 22
0 30 94 108
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U17B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
4498 0 0
2
5.90066e-315 5.46818e-315
0
9 2-In AND~
219 975 941 0 3 22
0 96 91 106
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
9728 0 0
2
5.90066e-315 5.47077e-315
0
9 2-In AND~
219 973 1037 0 3 22
0 32 93 104
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3789 0 0
2
5.90066e-315 5.47207e-315
0
8 3-In OR~
219 1070 980 0 4 22
0 106 105 104 98
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U2C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 12 0
1 U
3978 0 0
2
5.90066e-315 5.47336e-315
0
9 2-In AND~
219 974 991 0 3 22
0 91 93 105
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3494 0 0
2
5.90066e-315 5.47466e-315
0
9 2-In AND~
219 972 1099 0 3 22
0 96 31 103
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
3507 0 0
2
5.90066e-315 5.47595e-315
0
9 2-In AND~
219 970 1195 0 3 22
0 32 92 101
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
5151 0 0
2
5.90066e-315 5.47725e-315
0
8 3-In OR~
219 1067 1138 0 4 22
0 103 102 101 97
0
0 0 608 0
4 4075
-14 -24 14 -16
4 U19A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 15 0
1 U
3701 0 0
2
5.90066e-315 5.47854e-315
0
9 2-In AND~
219 971 1149 0 3 22
0 31 92 102
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
8585 0 0
2
5.90066e-315 5.47984e-315
0
9 Inverter~
13 499 1227 0 2 22
0 32 96
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U14F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
8809 0 0
2
5.90066e-315 5.48113e-315
0
9 Inverter~
13 1854 735 0 2 22
0 69 85
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U20A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 16 0
1 U
5993 0 0
2
5.90066e-315 5.48243e-315
0
14 Logic Display~
6 2088 681 0 1 2
10 79
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8654 0 0
2
5.90066e-315 5.48372e-315
0
14 Logic Display~
6 2358 681 0 1 2
10 73
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7223 0 0
2
5.90066e-315 5.48502e-315
0
14 Logic Display~
6 2393 680 0 1 2
10 72
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
5.90066e-315 5.48631e-315
0
14 Logic Display~
6 2425 680 0 1 2
10 71
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3104 0 0
2
5.90066e-315 5.48761e-315
0
14 Logic Display~
6 2458 681 0 1 2
10 70
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3296 0 0
2
5.90066e-315 5.4889e-315
0
14 Logic Display~
6 2189 681 0 1 2
10 77
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
5.90066e-315 5.4902e-315
0
14 Logic Display~
6 2224 680 0 1 2
10 76
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
949 0 0
2
5.90066e-315 5.49149e-315
0
14 Logic Display~
6 2256 680 0 1 2
10 75
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3371 0 0
2
5.90066e-315 5.49279e-315
0
14 Logic Display~
6 2289 681 0 1 2
10 74
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7311 0 0
2
5.90066e-315 5.49408e-315
0
14 Logic Display~
6 2021 682 0 1 2
10 81
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90066e-315 5.49538e-315
0
14 Logic Display~
6 2056 681 0 1 2
10 80
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3526 0 0
2
5.90066e-315 5.49667e-315
0
14 Logic Display~
6 2121 682 0 1 2
10 78
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4129 0 0
2
5.90066e-315 5.49797e-315
0
14 Logic Display~
6 1957 684 0 1 2
10 82
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6278 0 0
2
5.90066e-315 5.49926e-315
0
14 Logic Display~
6 1924 683 0 1 2
10 83
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
5.90066e-315 5.50056e-315
0
14 Logic Display~
6 1892 683 0 1 2
10 84
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8323 0 0
2
5.90066e-315 5.50185e-315
0
14 Logic Display~
6 1857 684 0 1 2
22 85
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-6 -19 8 -11
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3984 0 0
2
5.90066e-315 5.50315e-315
0
9 Inverter~
13 1889 731 0 2 22
0 68 84
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U20B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 16 0
1 U
7622 0 0
2
5.90066e-315 5.50444e-315
0
9 Inverter~
13 1921 732 0 2 22
0 67 83
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U20C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 16 0
1 U
816 0 0
2
5.90066e-315 5.50574e-315
0
9 Inverter~
13 1954 731 0 2 22
0 66 82
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U20D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 16 0
1 U
4656 0 0
2
5.90066e-315 5.50703e-315
0
9 Inverter~
13 2118 727 0 2 22
0 62 78
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U20E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 16 0
1 U
6356 0 0
2
5.90066e-315 5.50833e-315
0
9 Inverter~
13 2085 728 0 2 22
0 63 79
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U20F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 16 0
1 U
7479 0 0
2
5.90066e-315 5.50963e-315
0
9 Inverter~
13 2053 727 0 2 22
0 64 80
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U21A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 17 0
1 U
5690 0 0
2
5.90066e-315 5.51092e-315
0
9 Inverter~
13 2018 731 0 2 22
0 65 81
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U21B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 17 0
1 U
5617 0 0
2
5.90066e-315 5.51222e-315
0
9 Inverter~
13 2287 726 0 2 22
0 58 74
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U21C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 17 0
1 U
3903 0 0
2
5.90066e-315 5.51286e-315
0
9 Inverter~
13 2254 727 0 2 22
0 59 75
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U21D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 17 0
1 U
4452 0 0
2
5.90066e-315 5.51351e-315
0
9 Inverter~
13 2222 726 0 2 22
0 60 76
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U21E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 17 0
1 U
6282 0 0
2
5.90066e-315 5.51416e-315
0
9 Inverter~
13 2187 730 0 2 22
0 61 77
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U21F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 17 0
1 U
7187 0 0
2
5.90066e-315 5.51481e-315
0
9 Inverter~
13 2456 726 0 2 22
0 54 70
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U22A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 18 0
1 U
6866 0 0
2
5.90066e-315 5.51545e-315
0
9 Inverter~
13 2423 727 0 2 22
0 55 71
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U22B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 18 0
1 U
7670 0 0
2
5.90066e-315 5.5161e-315
0
9 Inverter~
13 2391 726 0 2 22
0 56 72
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U22C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 18 0
1 U
951 0 0
2
5.90066e-315 5.51675e-315
0
9 Inverter~
13 2356 730 0 2 22
0 57 73
0
0 0 96 90
6 74LS04
-21 -19 21 -11
4 U22D
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 18 0
1 U
9536 0 0
2
5.90066e-315 5.5174e-315
0
7 Pulser~
4 1122 891 0 10 12
0 119 120 29 121 0 0 5 5 6
7
0
0 0 4640 0
0
3 V19
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5495 0 0
2
5.90066e-315 5.51804e-315
0
7 Ground~
168 603 421 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8152 0 0
2
5.90066e-315 5.51869e-315
0
8 2-In OR~
219 580 136 0 3 22
0 13 25 51
0
0 0 96 270
6 74LS32
-21 -24 21 -16
4 U12B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6223 0 0
2
5.90066e-315 5.51934e-315
0
8 2-In OR~
219 642 134 0 3 22
0 12 24 50
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U12C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
5441 0 0
2
5.90066e-315 5.51999e-315
0
8 2-In OR~
219 723 134 0 3 22
0 11 23 49
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U12D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3189 0 0
2
5.90066e-315 5.52063e-315
0
8 2-In OR~
219 786 132 0 3 22
0 10 22 48
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U13A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8460 0 0
2
5.90066e-315 5.52128e-315
0
8 2-In OR~
219 869 130 0 3 22
0 6 20 47
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U13B
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
5179 0 0
2
5.90066e-315 5.52193e-315
0
8 2-In OR~
219 926 130 0 3 22
0 5 19 46
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U13C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3593 0 0
2
5.90066e-315 5.52258e-315
0
8 2-In OR~
219 1010 131 0 3 22
0 4 18 45
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U13D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3928 0 0
2
5.90066e-315 5.52322e-315
0
8 2-In OR~
219 1075 134 0 3 22
0 3 17 44
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U15A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
363 0 0
2
5.90066e-315 5.52387e-315
0
9 Inverter~
13 583 221 0 2 22
0 51 43
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U22E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 18 0
1 U
8132 0 0
2
5.90066e-315 5.52452e-315
0
9 Inverter~
13 640 220 0 2 22
0 50 42
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U22F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 18 0
1 U
65 0 0
2
5.90066e-315 5.52517e-315
0
9 Inverter~
13 724 222 0 2 22
0 49 41
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U16A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
6609 0 0
2
5.90066e-315 5.52581e-315
0
9 Inverter~
13 785 221 0 2 22
0 48 40
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U23A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 19 0
1 U
8995 0 0
2
5.90066e-315 5.52646e-315
0
9 Inverter~
13 867 221 0 2 22
0 47 39
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U23B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 19 0
1 U
3918 0 0
2
5.90066e-315 5.52711e-315
0
9 Inverter~
13 930 222 0 2 22
0 46 38
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U23C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 19 0
1 U
7519 0 0
2
5.90066e-315 5.52776e-315
0
9 Inverter~
13 1010 222 0 2 22
0 45 37
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U23D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 19 0
1 U
377 0 0
2
5.90066e-315 5.52841e-315
0
9 Inverter~
13 1075 221 0 2 22
0 44 36
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U23E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 19 0
1 U
8816 0 0
2
5.90066e-315 5.52905e-315
0
7 Ground~
168 804 386 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3877 0 0
2
5.90066e-315 5.5297e-315
0
9 2-In AND~
219 1204 893 0 3 22
0 26 29 28
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U24A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
926 0 0
2
5.90066e-315 5.53035e-315
0
9 Inverter~
13 825 461 0 2 22
0 27 26
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U23F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 19 0
1 U
7262 0 0
2
5.90066e-315 5.531e-315
0
9 Resistor~
219 1878 162 0 4 5
0 6 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R24
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5267 0 0
2
44974.8 18
0
9 Resistor~
219 1879 267 0 2 5
0 5 8
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R23
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8838 0 0
2
44974.8 19
0
9 Resistor~
219 1880 373 0 2 5
0 4 9
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R22
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7159 0 0
2
44974.8 20
0
9 Resistor~
219 2007 503 0 3 5
0 2 3 -1
0
0 0 864 90
2 1k
11 0 25 8
3 R21
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5812 0 0
2
44974.8 21
0
9 Resistor~
219 1631 164 0 4 5
0 13 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R20
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
331 0 0
2
44974.8 22
0
9 Resistor~
219 1632 269 0 2 5
0 12 15
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R19
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9604 0 0
2
44974.8 23
0
9 Resistor~
219 1633 375 0 2 5
0 11 16
0
0 0 864 180
2 1k
-7 -14 7 -6
3 R18
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7518 0 0
2
44974.8 24
0
9 Resistor~
219 1760 505 0 3 5
0 2 10 -1
0
0 0 864 90
2 1k
11 0 25 8
3 R17
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4832 0 0
2
44974.8 25
0
9 Resistor~
219 208 1179 0 3 5
0 2 17 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6798 0 0
2
44974.8 26
0
9 Resistor~
219 81 1049 0 4 5
0 18 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3336 0 0
2
44974.8 27
0
9 Resistor~
219 80 943 0 4 5
0 19 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8370 0 0
2
44974.8 28
0
9 Resistor~
219 79 838 0 4 5
0 20 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3910 0 0
2
44974.8 29
0
9 Resistor~
219 89 150 0 4 5
0 25 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
316 0 0
2
5.90066e-315 5.53164e-315
0
9 Resistor~
219 90 255 0 4 5
0 24 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
536 0 0
2
5.90066e-315 5.53229e-315
0
9 Resistor~
219 91 361 0 4 5
0 23 2 0 -1
0
0 0 864 180
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4460 0 0
2
5.90066e-315 5.53294e-315
0
9 Resistor~
219 218 491 0 3 5
0 2 22 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3260 0 0
2
5.90066e-315 5.53359e-315
0
193
0 4 3 0 0 8192 0 0 37 10 0 7
1994 452
1994 257
1255 257
1255 266
1163 266
1163 255
1196 255
0 3 4 0 0 8192 0 0 37 12 0 5
1940 373
1940 362
1168 362
1168 246
1196 246
0 2 5 0 0 8192 0 0 37 8 0 7
1947 267
1947 257
1250 257
1250 261
1173 261
1173 237
1196 237
0 1 6 0 0 8192 0 0 37 17 0 5
1946 162
1946 221
1173 221
1173 228
1196 228
0 1 3 0 0 12416 0 0 101 10 0 5
2007 452
2001 452
2001 103
1087 103
1087 118
0 1 5 0 0 8320 0 0 99 8 0 4
1986 247
1986 99
938 99
938 114
0 1 6 0 0 12416 0 0 98 17 0 5
1989 143
1985 143
1985 94
881 94
881 114
1 1 5 0 0 0 0 114 9 0 0 4
1897 267
1986 267
1986 247
1978 247
0 2 7 0 0 4096 0 0 9 21 0 2
1822 247
1944 247
2 1 3 0 0 0 0 116 10 0 0 3
2007 485
2007 452
1980 452
0 2 7 0 0 4112 0 0 10 21 0 3
1822 450
1946 450
1946 452
1 1 4 0 0 0 0 11 115 0 0 4
1977 352
1981 352
1981 373
1898 373
0 2 7 0 0 0 0 0 11 21 0 2
1822 352
1943 352
1 1 4 0 0 8320 0 100 11 0 0 5
1022 115
1022 95
1995 95
1995 352
1977 352
1 2 2 0 0 12288 0 12 113 0 0 5
2007 549
2007 525
1847 525
1847 162
1860 162
1 1 2 0 0 0 0 12 116 0 0 2
2007 549
2007 521
1 1 6 0 0 0 0 113 13 0 0 4
1896 162
1989 162
1989 142
1981 142
0 2 7 0 0 4096 0 0 13 21 0 2
1822 142
1947 142
0 2 8 0 0 4224 0 0 114 0 0 2
1851 267
1861 267
0 2 9 0 0 4224 0 0 115 0 0 2
1851 373
1862 373
1 0 7 0 0 4224 0 8 0 0 0 2
1822 87
1822 737
4 0 10 0 0 12288 0 36 0 0 31 4
1194 176
1180 176
1180 479
1760 479
3 0 11 0 0 12288 0 36 0 0 33 5
1194 167
1185 167
1185 384
1693 384
1693 375
2 0 12 0 0 12288 0 36 0 0 29 5
1194 158
1190 158
1190 278
1696 278
1696 269
1 0 13 0 0 12288 0 36 0 0 38 5
1194 149
1190 149
1190 122
1695 122
1695 164
0 1 10 0 0 12416 0 0 97 31 0 5
1760 456
1754 456
1754 96
798 96
798 116
0 1 12 0 0 8320 0 0 95 29 0 4
1739 249
1739 93
654 93
654 118
0 1 13 0 0 12416 0 0 94 38 0 5
1742 146
1738 146
1738 93
592 93
592 120
1 1 12 0 0 0 0 118 15 0 0 4
1650 269
1739 269
1739 249
1731 249
0 2 14 0 0 4096 0 0 15 42 0 2
1575 249
1697 249
2 1 10 0 0 0 0 120 16 0 0 3
1760 487
1760 454
1733 454
0 2 14 0 0 4096 0 0 16 42 0 2
1575 454
1699 454
1 1 11 0 0 0 0 17 119 0 0 4
1730 354
1734 354
1734 375
1651 375
0 2 14 0 0 0 0 0 17 42 0 2
1575 354
1696 354
1 1 11 0 0 8320 0 96 17 0 0 5
735 118
735 93
1748 93
1748 354
1730 354
1 2 2 0 0 0 0 18 117 0 0 5
1760 551
1760 527
1600 527
1600 164
1613 164
1 1 2 0 0 0 0 18 120 0 0 2
1760 551
1760 523
1 1 13 0 0 0 0 117 19 0 0 4
1649 164
1742 164
1742 144
1734 144
0 2 14 0 0 4096 0 0 19 42 0 2
1575 144
1700 144
0 2 15 0 0 4224 0 0 118 0 0 2
1604 269
1614 269
0 2 16 0 0 4224 0 0 119 0 0 2
1604 375
1615 375
1 0 14 0 0 4224 0 14 0 0 0 2
1575 89
1575 739
2 0 17 0 0 12416 0 101 0 0 59 5
1069 118
1069 47
342 47
342 1128
208 1128
2 0 18 0 0 12416 0 100 0 0 53 6
1004 115
1004 87
197 87
197 1023
192 1023
192 1028
0 2 19 0 0 8320 0 0 99 56 0 5
193 923
911 923
911 99
920 99
920 114
0 2 20 0 0 8320 0 0 98 54 0 5
194 820
855 820
855 99
863 99
863 114
1 1 18 0 0 0 0 22 122 0 0 4
178 1028
182 1028
182 1049
99 1049
2 0 21 0 0 4096 0 23 0 0 52 2
147 1128
25 1128
2 0 21 0 0 0 0 22 0 0 52 2
144 1028
25 1028
2 0 21 0 0 4096 0 20 0 0 52 2
148 818
25 818
2 0 21 0 0 0 0 24 0 0 52 2
145 923
25 923
0 0 21 0 0 8192 0 0 0 70 0 3
27 763
25 763
25 1413
1 0 18 0 0 0 0 22 0 0 0 2
178 1028
196 1028
1 1 20 0 0 0 0 124 20 0 0 4
97 838
194 838
194 818
182 818
2 1 2 0 0 8320 0 124 21 0 0 5
61 838
52 838
52 1216
208 1216
208 1225
1 1 19 0 0 0 0 123 24 0 0 4
98 943
193 943
193 923
179 923
2 0 2 0 0 0 0 123 0 0 55 2
62 943
52 943
2 0 2 0 0 0 0 122 0 0 55 2
63 1049
52 1049
2 1 17 0 0 0 0 121 23 0 0 3
208 1161
208 1128
181 1128
1 1 2 0 0 0 0 21 121 0 0 2
208 1225
208 1197
0 2 22 0 0 4224 0 0 97 77 0 5
218 441
773 441
773 101
780 101
780 116
0 2 23 0 0 8320 0 0 96 71 0 4
201 340
201 93
717 93
717 118
0 2 24 0 0 4224 0 0 95 74 0 5
203 235
565 235
565 98
636 98
636 118
0 2 25 0 0 4224 0 0 94 72 0 5
204 130
571 130
571 105
574 105
574 120
1 1 23 0 0 0 0 28 127 0 0 4
188 340
192 340
192 361
109 361
2 0 21 0 0 0 0 27 0 0 70 2
157 440
27 440
2 0 21 0 0 0 0 28 0 0 70 2
154 340
27 340
2 0 21 0 0 0 0 30 0 0 70 2
158 130
27 130
2 0 21 0 0 0 0 26 0 0 70 2
155 235
27 235
1 0 21 0 0 8320 0 25 0 0 52 4
33 75
27 75
27 768
25 768
1 0 23 0 0 0 0 28 0 0 0 2
188 340
206 340
1 1 25 0 0 0 0 125 30 0 0 4
107 150
204 150
204 130
192 130
2 1 2 0 0 0 0 125 29 0 0 5
71 150
62 150
62 528
218 528
218 537
1 1 24 0 0 0 0 126 26 0 0 4
108 255
203 255
203 235
189 235
2 0 2 0 0 0 0 126 0 0 73 2
72 255
62 255
2 0 2 0 0 0 0 127 0 0 73 2
73 361
62 361
2 1 22 0 0 0 0 128 27 0 0 3
218 473
218 440
191 440
1 1 2 0 0 0 0 29 128 0 0 2
218 537
218 509
2 1 26 0 0 8320 0 112 111 0 0 6
846 461
1153 461
1153 869
1167 869
1167 884
1180 884
14 1 27 0 0 8320 0 31 112 0 0 3
732 428
732 461
810 461
3 2 28 0 0 8320 0 111 40 0 0 6
1225 893
1239 893
1239 1171
1156 1171
1156 1156
1164 1156
3 2 28 0 0 0 0 111 39 0 0 6
1225 893
1234 893
1234 1013
1154 1013
1154 998
1162 998
0 2 28 0 0 0 0 0 42 84 0 5
1229 893
1229 689
1150 689
1150 674
1158 674
3 2 28 0 0 0 0 111 41 0 0 6
1225 893
1229 893
1229 846
1146 846
1146 831
1159 831
3 2 29 0 0 4224 0 92 111 0 0 4
1146 882
1172 882
1172 902
1180 902
1 0 30 0 0 4096 0 50 0 0 87 3
949 816
900 816
900 784
2 2 30 0 0 4224 0 35 47 0 0 3
727 512
727 784
950 784
1 0 31 0 0 4096 0 58 0 0 89 3
947 1140
910 1140
910 1108
2 2 31 0 0 4224 0 33 55 0 0 3
665 511
665 1108
948 1108
1 0 32 0 0 4096 0 56 0 0 191 2
946 1186
529 1186
1 0 32 0 0 4096 0 52 0 0 191 2
949 1028
529 1028
1 0 32 0 0 0 0 48 0 0 191 2
948 862
529 862
1 0 32 0 0 4096 0 45 0 0 191 2
950 701
529 701
1 1 2 0 0 0 0 31 110 0 0 4
732 352
732 348
804 348
804 380
13 1 33 0 0 4224 0 31 35 0 0 4
705 428
705 468
727 468
727 476
12 1 34 0 0 4224 0 31 34 0 0 2
696 428
696 476
11 1 35 0 0 4224 0 31 33 0 0 4
687 428
687 467
665 467
665 475
2 2 36 0 0 8320 0 109 31 0 0 4
1078 239
1078 320
714 320
714 352
2 3 37 0 0 8320 0 108 31 0 0 4
1013 240
1013 325
705 325
705 352
2 4 38 0 0 8320 0 107 31 0 0 4
933 240
933 330
696 330
696 352
2 5 39 0 0 8320 0 106 31 0 0 4
870 239
870 335
687 335
687 352
2 6 40 0 0 8320 0 105 31 0 0 4
788 239
788 339
678 339
678 352
2 7 41 0 0 4224 0 104 31 0 0 4
727 240
727 344
669 344
669 352
2 8 42 0 0 4224 0 103 31 0 0 4
643 238
643 339
660 339
660 352
2 9 43 0 0 4224 0 102 31 0 0 4
586 239
586 344
651 344
651 352
3 1 44 0 0 4224 0 101 109 0 0 2
1078 164
1078 203
3 1 45 0 0 4224 0 100 108 0 0 2
1013 161
1013 204
3 1 46 0 0 4224 0 99 107 0 0 4
929 160
929 196
933 196
933 204
3 1 47 0 0 4224 0 98 106 0 0 4
872 160
872 195
870 195
870 203
3 1 48 0 0 4224 0 97 105 0 0 4
789 162
789 195
788 195
788 203
3 1 49 0 0 4224 0 96 104 0 0 4
726 164
726 196
727 196
727 204
3 1 50 0 0 4224 0 95 103 0 0 4
645 164
645 194
643 194
643 202
3 1 51 0 0 4224 0 94 102 0 0 4
583 166
583 195
586 195
586 203
10 1 2 0 0 0 0 31 93 0 0 6
651 428
651 436
620 436
620 401
603 401
603 415
1 2 52 0 0 8320 0 7 32 0 0 4
1468 874
1498 874
1498 920
1540 920
1 1 53 0 0 8320 0 6 32 0 0 4
1468 837
1511 837
1511 911
1540 911
7 1 54 0 0 4224 0 32 88 0 0 3
1616 866
2459 866
2459 744
8 1 55 0 0 4224 0 32 89 0 0 3
1616 875
2426 875
2426 745
9 1 56 0 0 4224 0 32 90 0 0 3
1616 884
2394 884
2394 744
10 1 57 0 0 4224 0 32 91 0 0 3
1616 893
2359 893
2359 748
11 1 58 0 0 4224 0 32 84 0 0 3
1616 902
2290 902
2290 744
12 1 59 0 0 4224 0 32 85 0 0 3
1616 911
2257 911
2257 745
13 1 60 0 0 4224 0 32 86 0 0 3
1616 920
2225 920
2225 744
14 1 61 0 0 4224 0 32 87 0 0 3
1616 929
2190 929
2190 748
15 1 62 0 0 4224 0 32 80 0 0 3
1616 938
2121 938
2121 745
16 1 63 0 0 4224 0 32 81 0 0 3
1616 947
2088 947
2088 746
17 1 64 0 0 4224 0 32 82 0 0 3
1616 956
2056 956
2056 745
18 1 65 0 0 4224 0 32 83 0 0 3
1616 965
2021 965
2021 749
19 1 66 0 0 4224 0 32 79 0 0 3
1616 974
1957 974
1957 749
20 1 67 0 0 4224 0 32 78 0 0 3
1616 983
1924 983
1924 750
21 1 68 0 0 4224 0 32 77 0 0 3
1616 992
1892 992
1892 749
22 1 69 0 0 8320 0 32 60 0 0 3
1616 1001
1857 1001
1857 753
1 2 70 0 0 8320 0 65 88 0 0 3
2458 699
2459 699
2459 708
1 2 71 0 0 8320 0 64 89 0 0 3
2425 698
2426 698
2426 709
1 2 72 0 0 8320 0 63 90 0 0 3
2393 698
2394 698
2394 708
1 2 73 0 0 8320 0 62 91 0 0 3
2358 699
2359 699
2359 712
1 2 74 0 0 8320 0 69 84 0 0 3
2289 699
2290 699
2290 708
1 2 75 0 0 8320 0 68 85 0 0 3
2256 698
2257 698
2257 709
1 2 76 0 0 8320 0 67 86 0 0 3
2224 698
2225 698
2225 708
1 2 77 0 0 8320 0 66 87 0 0 3
2189 699
2190 699
2190 712
1 2 78 0 0 4224 0 72 80 0 0 2
2121 700
2121 709
1 2 79 0 0 4224 0 61 81 0 0 2
2088 699
2088 710
1 2 80 0 0 4224 0 71 82 0 0 2
2056 699
2056 709
1 2 81 0 0 4224 0 70 83 0 0 2
2021 700
2021 713
1 2 82 0 0 4224 0 73 79 0 0 2
1957 702
1957 713
1 2 83 0 0 4224 0 74 78 0 0 2
1924 701
1924 714
1 2 84 0 0 4224 0 75 77 0 0 2
1892 701
1892 713
1 2 85 0 0 4224 0 76 60 0 0 2
1857 702
1857 717
4 6 86 0 0 4224 0 40 32 0 0 4
1212 1138
1389 1138
1389 974
1546 974
4 5 87 0 0 12416 0 39 32 0 0 4
1210 980
1366 980
1366 965
1546 965
4 4 88 0 0 12416 0 41 32 0 0 4
1207 813
1365 813
1365 956
1546 956
4 3 89 0 0 8320 0 42 32 0 0 4
1206 656
1389 656
1389 947
1546 947
1 0 90 0 0 8192 0 43 0 0 164 3
951 655
929 655
929 623
1 0 91 0 0 4096 0 54 0 0 155 3
950 982
910 982
910 950
2 2 91 0 0 4224 0 34 51 0 0 3
696 512
696 950
951 950
2 0 92 0 0 4096 0 56 0 0 187 2
946 1204
788 1204
2 0 92 0 0 4096 0 58 0 0 187 2
947 1158
788 1158
2 0 93 0 0 4096 0 52 0 0 188 2
949 1046
717 1046
2 0 93 0 0 4096 0 54 0 0 188 2
950 1000
717 1000
2 0 94 0 0 4096 0 48 0 0 189 2
948 880
654 880
2 0 94 0 0 4096 0 50 0 0 189 2
949 834
654 834
2 0 95 0 0 4096 0 45 0 0 190 2
950 719
592 719
2 0 95 0 0 4096 0 43 0 0 190 2
951 673
592 673
3 2 90 0 0 12416 0 38 46 0 0 6
1327 201
1404 201
1404 447
914 447
914 623
952 623
1 0 96 0 0 4096 0 55 0 0 169 2
948 1090
502 1090
1 0 96 0 0 4096 0 51 0 0 169 2
951 932
502 932
1 0 96 0 0 0 0 47 0 0 169 2
950 766
502 766
1 0 96 0 0 4096 0 46 0 0 169 2
952 605
502 605
2 0 96 0 0 4224 0 59 0 0 0 2
502 1209
502 511
1 1 32 0 0 0 0 5 59 0 0 3
529 1259
502 1259
502 1245
4 1 97 0 0 4224 0 57 40 0 0 2
1100 1138
1164 1138
4 1 98 0 0 4224 0 53 39 0 0 2
1103 980
1162 980
4 1 99 0 0 8320 0 49 41 0 0 3
1102 814
1102 813
1159 813
4 1 100 0 0 8320 0 44 42 0 0 3
1104 653
1104 656
1158 656
3 3 101 0 0 4224 0 56 57 0 0 4
991 1195
1048 1195
1048 1147
1054 1147
3 2 102 0 0 4224 0 58 57 0 0 4
992 1149
1036 1149
1036 1138
1055 1138
3 1 103 0 0 4224 0 55 57 0 0 4
993 1099
1031 1099
1031 1129
1054 1129
3 3 104 0 0 4224 0 52 53 0 0 4
994 1037
1051 1037
1051 989
1057 989
3 2 105 0 0 4224 0 54 53 0 0 4
995 991
1039 991
1039 980
1058 980
3 1 106 0 0 4224 0 51 53 0 0 4
996 941
1034 941
1034 971
1057 971
3 3 107 0 0 4224 0 48 49 0 0 4
993 871
1050 871
1050 823
1056 823
3 2 108 0 0 4224 0 50 49 0 0 4
994 825
1038 825
1038 814
1057 814
3 1 109 0 0 4224 0 47 49 0 0 4
995 775
1033 775
1033 805
1056 805
3 3 110 0 0 4224 0 45 44 0 0 4
995 710
1052 710
1052 662
1058 662
3 2 111 0 0 4224 0 43 44 0 0 4
996 664
1040 664
1040 653
1059 653
3 1 112 0 0 4224 0 46 44 0 0 4
997 614
1035 614
1035 644
1058 644
1 0 92 0 0 4224 0 1 0 0 0 2
788 1261
788 592
1 0 93 0 0 4224 0 2 0 0 0 2
717 1259
717 592
1 0 94 0 0 4224 0 3 0 0 0 2
654 1259
654 591
1 0 95 0 0 4224 0 4 0 0 0 2
592 1262
592 509
1 0 32 0 0 4224 0 5 0 0 0 2
529 1259
529 509
5 2 113 0 0 8320 0 37 38 0 0 4
1246 241
1257 241
1257 210
1281 210
5 1 114 0 0 8320 0 36 38 0 0 4
1244 162
1257 162
1257 192
1281 192
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
