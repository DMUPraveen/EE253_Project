CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 10 30 100 10
2 80 1278 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
170 176 283 273
9437202 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 861 129 0 1 11
0 4
0
0 0 20848 270
2 0V
-6 -21 8 -13
2 V1
11 -15 25 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9730 0 0
2
44971.9 1
0
13 Logic Switch~
5 111 154 0 1 11
0 20
0
0 0 20848 90
2 0V
11 -5 25 3
3 V16
8 -15 29 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9874 0 0
2
5.90066e-315 5.37752e-315
0
13 Logic Switch~
5 152 154 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 20848 90
2 5V
11 -5 25 3
3 V15
8 -15 29 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
364 0 0
2
5.90066e-315 5.36716e-315
0
13 Logic Switch~
5 196 155 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 20848 90
2 5V
11 -5 25 3
3 V14
8 -15 29 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3656 0 0
2
5.90066e-315 5.3568e-315
0
13 Logic Switch~
5 236 155 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 20848 90
2 5V
11 -5 25 3
3 V13
8 -15 29 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3131 0 0
2
5.90066e-315 5.34643e-315
0
13 Logic Switch~
5 315 154 0 1 11
0 19
0
0 0 20848 90
2 0V
11 -5 25 3
3 V12
8 -15 29 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6772 0 0
2
5.90066e-315 5.32571e-315
0
13 Logic Switch~
5 359 155 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 20848 90
2 5V
11 -5 25 3
3 V11
8 -15 29 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9557 0 0
2
5.90066e-315 5.30499e-315
0
13 Logic Switch~
5 401 155 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 20848 90
2 5V
11 -5 25 3
3 V10
8 -15 29 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5789 0 0
2
5.90066e-315 5.26354e-315
0
13 Logic Switch~
5 445 156 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 20848 90
2 5V
11 -5 25 3
2 V9
11 -15 25 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7328 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 951 361 0 1 2
14 2
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 R3
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4799 0 0
2
44971.9 0
0
14 Logic Display~
6 956 191 0 1 2
10 3
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 R1
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9196 0 0
2
44971.9 0
0
14 Logic Display~
6 861 61 0 1 2
22 4
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 R2
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3857 0 0
2
44971.9 0
0
9 2-In AND~
219 869 365 0 3 22
0 4 6 2
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 A28
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7125 0 0
2
5.90066e-315 0
0
9 2-In AND~
219 868 196 0 3 22
0 4 5 3
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 A29
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3641 0 0
2
5.90066e-315 0
0
9 Inverter~
13 787 244 0 2 22
0 6 5
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 A30
-11 -29 10 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9821 0 0
2
5.90066e-315 0
0
8 2-In OR~
219 674 302 0 3 22
0 8 7 6
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 A31
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3187 0 0
2
5.90066e-315 0
0
8 2-In OR~
219 589 360 0 3 22
0 10 9 7
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 A32
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
762 0 0
2
5.90066e-315 0
0
8 2-In OR~
219 594 244 0 3 22
0 12 11 8
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 A33
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
39 0 0
2
5.90066e-315 0
0
6 74136~
219 501 402 0 3 22
0 14 13 9
0
0 0 112 0
7 74LS136
-24 -24 25 -16
3 A34
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9450 0 0
2
5.90066e-315 0
0
6 74136~
219 498 337 0 3 22
0 16 15 10
0
0 0 112 0
7 74LS136
-24 -24 25 -16
3 A35
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3236 0 0
2
5.90066e-315 0
0
6 74136~
219 498 273 0 3 22
0 18 17 11
0
0 0 112 0
7 74LS136
-24 -24 25 -16
3 A36
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3321 0 0
2
5.90066e-315 0
0
6 74136~
219 499 211 0 3 22
0 20 19 12
0
0 0 112 0
7 74LS136
-24 -24 25 -16
3 A37
-10 -34 11 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8879 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 112 97 0 1 2
15 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5433 0 0
2
5.90066e-315 5.42414e-315
0
14 Logic Display~
6 153 97 0 1 2
15 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3679 0 0
2
5.90066e-315 5.41896e-315
0
14 Logic Display~
6 197 98 0 1 2
15 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9342 0 0
2
5.90066e-315 5.41378e-315
0
14 Logic Display~
6 237 98 0 1 2
15 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 N0
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3623 0 0
2
5.90066e-315 5.4086e-315
0
14 Logic Display~
6 316 97 0 1 2
12 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3722 0 0
2
5.90066e-315 5.40342e-315
0
14 Logic Display~
6 360 98 0 1 2
12 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8993 0 0
2
5.90066e-315 5.39824e-315
0
14 Logic Display~
6 402 98 0 1 2
12 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3723 0 0
2
5.90066e-315 5.39306e-315
0
14 Logic Display~
6 446 99 0 1 2
12 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6244 0 0
2
5.90066e-315 5.38788e-315
0
46
3 1 2 0 0 8320 0 13 10 0 0 5
890 365
904 365
904 412
951 412
951 379
3 1 3 0 0 8320 0 14 11 0 0 5
889 196
904 196
904 256
956 256
956 209
0 1 4 0 0 4224 0 0 13 4 0 3
830 141
830 356
845 356
1 1 4 0 0 0 0 1 14 0 0 4
861 141
807 141
807 187
844 187
1 1 4 0 0 0 0 12 1 0 0 4
861 79
903 79
903 141
861 141
2 2 5 0 0 4224 0 15 14 0 0 3
808 244
808 205
844 205
3 2 6 0 0 8320 0 16 13 0 0 3
707 302
707 374
845 374
3 1 6 0 0 0 0 16 15 0 0 3
707 302
707 244
772 244
3 2 7 0 0 4224 0 17 16 0 0 3
622 360
622 311
661 311
3 1 8 0 0 4224 0 18 16 0 0 3
627 244
627 293
661 293
3 2 9 0 0 8320 0 19 17 0 0 3
534 402
534 369
576 369
3 1 10 0 0 8320 0 20 17 0 0 3
531 337
531 351
576 351
3 2 11 0 0 8320 0 21 18 0 0 3
531 273
531 253
581 253
3 1 12 0 0 8320 0 22 18 0 0 3
532 211
532 235
581 235
2 0 13 0 0 4096 0 19 0 0 23 2
485 411
425 411
1 0 14 0 0 4096 0 19 0 0 27 2
485 393
215 393
2 0 15 0 0 4096 0 20 0 0 24 2
482 346
380 346
1 0 16 0 0 4096 0 20 0 0 28 2
482 328
174 328
2 0 17 0 0 4096 0 21 0 0 25 2
482 282
342 282
1 0 18 0 0 4096 0 21 0 0 29 2
482 264
135 264
2 0 19 0 0 4096 0 22 0 0 26 2
483 220
291 220
1 0 20 0 0 4096 0 22 0 0 30 2
483 202
93 202
0 0 13 0 0 8320 0 0 0 31 0 3
446 139
425 139
425 545
0 0 15 0 0 8320 0 0 0 33 0 3
402 137
380 137
380 542
0 0 17 0 0 8320 0 0 0 35 0 3
360 138
342 138
342 547
0 0 19 0 0 8320 0 0 0 37 0 3
316 136
291 136
291 544
0 0 14 0 0 8320 0 0 0 39 0 3
237 137
215 137
215 548
0 0 16 0 0 8320 0 0 0 41 0 3
197 138
174 138
174 546
0 0 18 0 0 8320 0 0 0 43 0 3
153 136
135 136
135 548
0 0 20 0 0 8320 0 0 0 45 0 3
112 137
93 137
93 547
1 0 13 0 0 0 0 30 0 0 32 2
446 117
446 139
1 1 13 0 0 0 0 9 30 0 0 2
446 143
446 117
1 0 15 0 0 0 0 29 0 0 34 2
402 116
402 138
1 1 15 0 0 0 0 8 29 0 0 2
402 142
402 116
1 0 17 0 0 0 0 28 0 0 36 2
360 116
360 138
1 1 17 0 0 0 0 7 28 0 0 2
360 142
360 116
1 0 19 0 0 0 0 27 0 0 38 2
316 115
316 137
1 1 19 0 0 0 0 6 27 0 0 2
316 141
316 115
1 0 14 0 0 0 0 26 0 0 40 2
237 116
237 138
1 1 14 0 0 0 0 5 26 0 0 2
237 142
237 116
1 0 16 0 0 0 0 25 0 0 42 2
197 116
197 138
1 1 16 0 0 0 0 4 25 0 0 2
197 142
197 116
1 0 18 0 0 0 0 24 0 0 44 2
153 115
153 137
1 1 18 0 0 0 0 3 24 0 0 2
153 141
153 115
1 0 20 0 0 0 0 23 0 0 46 2
112 115
112 137
1 1 20 0 0 0 0 2 23 0 0 2
112 141
112 115
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
984 363 1061 387
994 371 1050 387
7 UNEQUAL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
988 191 1049 215
998 199 1038 215
5 N = M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
869 43 916 67
880 52 904 68
4 USER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
369 47 394 71
377 55 385 71
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
163 50 188 74
171 58 179 74
1 N
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
118 26 235 50
128 34 224 50
12 FIRST NUMBER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
329 25 454 49
339 33 443 49
13 SECOND NUMBER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
