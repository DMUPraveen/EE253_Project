CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 0 30 130 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
23
12 SPST Switch~
165 372 42 0 2 11
0 4 5
0
0 0 4720 0
0
2 S5
-7 -18 7 -10
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
523 0 0
2
5.90066e-315 0
0
10 2-In NAND~
219 469 40 0 3 22
0 4 4 3
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6748 0 0
2
5.90066e-315 0
0
7 74LS245
64 536 104 0 18 37
0 23 24 25 26 27 28 29 30 31
32 33 34 6 7 8 9 3 35
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
6901 0 0
2
5.90066e-315 0
0
7 74LS245
64 523 322 0 18 37
0 36 37 38 39 10 11 12 13 40
41 42 43 6 7 8 9 4 5
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
842 0 0
2
5.90066e-315 0
0
7 Pulser~
4 528 451 0 10 12
0 44 45 14 46 0 0 5 5 6
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 1 0 0
1 V
3277 0 0
2
5.90066e-315 0
0
12 Quad D Flop~
47 667 217 0 9 19
0 9 8 7 6 18 17 16 15 14
0
0 0 4720 0
4 QDFF
-14 -44 14 -36
2 U4
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4212 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 788 151 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 763 151 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 734 151 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 706 151 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
5.90066e-315 0
0
6 74LS73
102 374 326 0 12 25
0 5 5 19 5 5 5 20 5 11
47 10 48
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
9592 0 0
2
5.90066e-315 0
0
6 74LS73
102 373 117 0 12 25
0 5 5 22 5 5 5 21 5 13
49 12 50
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
8748 0 0
2
5.90066e-315 0
0
14 NO PushButton~
191 171 207 0 2 5
0 21 5
0
0 0 4720 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7168 0 0
2
5.90066e-315 0
0
14 NO PushButton~
191 173 412 0 2 5
0 20 5
0
0 0 4720 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
631 0 0
2
5.90066e-315 0
0
14 NO PushButton~
191 170 312 0 2 5
0 19 5
0
0 0 4720 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9466 0 0
2
5.90066e-315 0
0
7 Ground~
168 217 523 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3266 0 0
2
5.90066e-315 0
0
14 NO PushButton~
191 174 102 0 2 5
0 22 5
0
0 0 4720 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7693 0 0
2
5.90066e-315 0
0
2 +V
167 266 26 0 1 3
0 5
0
0 0 54256 0
3 15V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3723 0 0
2
5.90066e-315 0
0
9 Resistor~
219 433 17 0 3 5
0 2 4 -1
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3440 0 0
2
5.90066e-315 0
0
9 Resistor~
219 88 130 0 4 5
0 22 2 0 -1
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6263 0 0
2
5.90066e-315 0
0
9 Resistor~
219 89 235 0 4 5
0 21 2 0 -1
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4900 0 0
2
5.90066e-315 0
0
9 Resistor~
219 90 341 0 4 5
0 19 2 0 -1
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8783 0 0
2
5.90066e-315 5.26354e-315
0
9 Resistor~
219 217 471 0 3 5
0 2 20 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3221 0 0
2
5.90066e-315 0
0
53
3 17 3 0 0 4224 0 2 3 0 0 3
496 40
496 68
498 68
0 17 4 0 0 4224 0 0 4 3 0 3
420 42
420 286
485 286
1 0 4 0 0 0 0 1 0 0 4 2
389 42
430 42
2 1 4 0 0 0 0 2 2 0 0 4
445 49
430 49
430 31
445 31
2 0 5 0 0 4096 0 1 0 0 52 3
355 42
267 42
267 46
1 0 2 0 0 12416 0 19 0 0 51 4
451 17
848 17
848 501
217 501
2 0 4 0 0 0 0 19 0 0 3 3
415 17
411 17
411 42
13 0 6 0 0 8320 0 3 0 0 12 3
568 113
571 113
571 227
14 0 7 0 0 8192 0 3 0 0 13 4
568 122
589 122
589 212
594 212
15 0 8 0 0 8192 0 3 0 0 14 4
568 131
608 131
608 199
613 199
16 0 9 0 0 4096 0 3 0 0 15 4
568 140
630 140
630 189
635 189
13 4 6 0 0 0 0 4 6 0 0 4
555 331
571 331
571 223
643 223
14 3 7 0 0 8320 0 4 6 0 0 4
555 340
594 340
594 211
643 211
15 2 8 0 0 8320 0 4 6 0 0 4
555 349
613 349
613 199
643 199
16 1 9 0 0 8320 0 4 6 0 0 4
555 358
635 358
635 187
643 187
11 5 10 0 0 12416 0 11 4 0 0 4
406 344
413 344
413 331
491 331
9 6 11 0 0 12416 0 11 4 0 0 4
406 308
425 308
425 340
491 340
11 7 12 0 0 8320 0 12 4 0 0 4
405 135
435 135
435 349
491 349
9 8 13 0 0 8320 0 12 4 0 0 4
405 99
449 99
449 358
491 358
3 9 14 0 0 8320 0 5 6 0 0 3
552 442
667 442
667 253
8 1 15 0 0 4224 0 6 7 0 0 3
691 223
788 223
788 169
7 1 16 0 0 4224 0 6 8 0 0 3
691 211
763 211
763 169
6 1 17 0 0 4224 0 6 9 0 0 3
691 199
734 199
734 169
5 1 18 0 0 8320 0 6 10 0 0 3
691 187
706 187
706 169
1 0 19 0 0 4096 0 15 0 0 45 2
187 320
205 320
8 0 5 0 0 0 0 11 0 0 53 4
336 362
265 362
265 360
267 360
7 1 20 0 0 12416 0 11 14 0 0 5
336 353
304 353
304 419
190 419
190 420
6 0 5 0 0 0 0 11 0 0 53 2
342 344
267 344
5 0 5 0 0 0 0 11 0 0 53 2
342 335
267 335
4 0 5 0 0 0 0 11 0 0 53 4
336 326
272 326
272 327
267 327
2 0 5 0 0 0 0 11 0 0 53 2
342 308
267 308
1 0 5 0 0 0 0 11 0 0 53 2
342 299
267 299
8 0 5 0 0 0 0 12 0 0 48 3
335 153
264 153
264 151
7 1 21 0 0 12416 0 12 13 0 0 4
335 144
303 144
303 215
188 215
6 0 5 0 0 0 0 12 0 0 53 2
341 135
267 135
5 0 5 0 0 0 0 12 0 0 53 2
341 126
267 126
4 0 5 0 0 0 0 12 0 0 53 4
335 117
271 117
271 118
267 118
3 0 22 0 0 4224 0 12 0 0 41 4
335 108
208 108
208 111
203 111
2 0 5 0 0 0 0 12 0 0 53 2
341 99
267 99
1 0 5 0 0 0 0 12 0 0 53 2
341 90
267 90
1 1 22 0 0 0 0 20 17 0 0 4
106 130
203 130
203 110
191 110
2 1 2 0 0 0 0 20 16 0 0 5
70 130
61 130
61 508
217 508
217 517
1 0 21 0 0 0 0 21 0 0 34 3
107 235
202 235
202 215
2 0 2 0 0 0 0 21 0 0 42 2
71 235
61 235
3 1 19 0 0 4224 0 11 22 0 0 6
336 317
209 317
209 320
205 320
205 341
108 341
2 0 2 0 0 0 0 22 0 0 42 2
72 341
61 341
2 0 20 0 0 0 0 23 0 0 27 2
217 453
217 419
2 0 5 0 0 12288 0 13 0 0 53 4
154 215
119 215
119 151
267 151
2 0 5 0 0 0 0 14 0 0 53 4
156 420
121 420
121 361
267 361
2 0 5 0 0 0 0 15 0 0 53 4
153 320
121 320
121 259
267 259
1 1 2 0 0 0 0 16 23 0 0 2
217 517
217 489
2 0 5 0 0 0 0 17 0 0 53 4
157 110
122 110
122 46
267 46
1 18 5 0 0 8320 0 18 4 0 0 6
266 35
267 35
267 405
559 405
559 286
555 286
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
